module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n906 , n907 , n908 , n909 , n910 , n911 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 ;
  assign n513 = ~x6 & ~x7 ;
  assign n514 = ~x5 & n513 ;
  assign n515 = ~x4 & n514 ;
  assign n516 = ~x3 & n515 ;
  assign n517 = ~x2 & n516 ;
  assign n518 = ~x1 & n517 ;
  assign n519 = ~x0 & n518 ;
  assign n520 = ~x15 & n519 ;
  assign n521 = ~x14 & n520 ;
  assign n522 = ~x13 & n521 ;
  assign n523 = ~x12 & n522 ;
  assign n524 = ~x11 & n523 ;
  assign n525 = ~x10 & n524 ;
  assign n526 = ~x9 & n525 ;
  assign n527 = ~x8 & n526 ;
  assign n528 = ~x23 & n527 ;
  assign n529 = ~x22 & n528 ;
  assign n530 = ~x21 & n529 ;
  assign n531 = ~x20 & n530 ;
  assign n532 = ~x19 & n531 ;
  assign n533 = ~x18 & n532 ;
  assign n534 = ~x17 & n533 ;
  assign n535 = ~x16 & n534 ;
  assign n536 = ~x31 & n535 ;
  assign n585 = n536 ^ x30 ;
  assign n541 = n534 ^ x16 ;
  assign n542 = n533 ^ x17 ;
  assign n543 = n532 ^ x18 ;
  assign n544 = n531 ^ x19 ;
  assign n545 = n530 ^ x20 ;
  assign n546 = n529 ^ x21 ;
  assign n547 = n528 ^ x22 ;
  assign n548 = n527 ^ x23 ;
  assign n549 = n526 ^ x8 ;
  assign n550 = n525 ^ x9 ;
  assign n551 = n523 ^ x11 ;
  assign n552 = n522 ^ x12 ;
  assign n553 = n521 ^ x13 ;
  assign n554 = n520 ^ x14 ;
  assign n555 = n519 ^ x15 ;
  assign n556 = n518 ^ x0 ;
  assign n557 = n517 ^ x1 ;
  assign n558 = n516 ^ x2 ;
  assign n559 = n514 ^ x4 ;
  assign n560 = n515 ^ x3 ;
  assign n561 = ~n559 & ~n560 ;
  assign n562 = ~n558 & n561 ;
  assign n563 = ~n557 & n562 ;
  assign n564 = n556 & ~n563 ;
  assign n565 = n555 & n564 ;
  assign n566 = n554 & n565 ;
  assign n567 = ~n553 & ~n566 ;
  assign n568 = n552 & ~n567 ;
  assign n569 = n551 & n568 ;
  assign n570 = n524 ^ x10 ;
  assign n571 = ~n569 & ~n570 ;
  assign n572 = n550 & ~n571 ;
  assign n573 = ~n549 & ~n572 ;
  assign n574 = n548 & ~n573 ;
  assign n575 = ~n547 & ~n574 ;
  assign n576 = n546 & ~n575 ;
  assign n577 = ~n545 & ~n576 ;
  assign n578 = n544 & ~n577 ;
  assign n579 = ~n543 & ~n578 ;
  assign n580 = ~n542 & n579 ;
  assign n581 = n535 ^ x31 ;
  assign n582 = ~n580 & ~n581 ;
  assign n583 = n541 & n582 ;
  assign n584 = n583 ^ n581 ;
  assign n592 = n585 ^ n584 ;
  assign n637 = n566 ^ n553 ;
  assign n619 = n565 ^ n554 ;
  assign n620 = n564 ^ n555 ;
  assign n621 = n563 ^ n556 ;
  assign n622 = n562 ^ n557 ;
  assign n623 = n561 ^ n558 ;
  assign n624 = n513 ^ x5 ;
  assign n586 = ~n584 & ~n585 ;
  assign n537 = ~x30 & n536 ;
  assign n587 = n537 ^ x29 ;
  assign n588 = n586 & ~n587 ;
  assign n538 = ~x29 & n537 ;
  assign n589 = n538 ^ x28 ;
  assign n590 = ~n588 & n589 ;
  assign n539 = ~x28 & n538 ;
  assign n540 = n539 ^ x27 ;
  assign n591 = n590 ^ n540 ;
  assign n593 = n587 ^ n586 ;
  assign n594 = ~n592 & n593 ;
  assign n595 = n589 ^ n588 ;
  assign n596 = n594 & ~n595 ;
  assign n597 = n591 & ~n596 ;
  assign n600 = ~n540 & ~n590 ;
  assign n598 = ~x27 & n539 ;
  assign n599 = n598 ^ x26 ;
  assign n601 = n600 ^ n599 ;
  assign n602 = ~n597 & ~n601 ;
  assign n604 = ~x26 & n598 ;
  assign n605 = n604 ^ x25 ;
  assign n603 = n599 & ~n600 ;
  assign n606 = n605 ^ n603 ;
  assign n607 = n602 & ~n606 ;
  assign n610 = x25 ^ x24 ;
  assign n608 = n604 ^ n603 ;
  assign n609 = ~n605 & n608 ;
  assign n611 = n610 ^ n609 ;
  assign n612 = n607 & ~n611 ;
  assign n625 = x7 & ~n612 ;
  assign n626 = ~x6 & n625 ;
  assign n627 = ~n624 & n626 ;
  assign n628 = n627 ^ n560 ;
  assign n629 = ~n559 & ~n628 ;
  assign n630 = n629 ^ n560 ;
  assign n631 = ~n561 & ~n630 ;
  assign n632 = n623 & ~n631 ;
  assign n633 = ~n622 & ~n632 ;
  assign n634 = ~n621 & ~n633 ;
  assign n635 = ~n620 & ~n634 ;
  assign n636 = ~n619 & n635 ;
  assign n651 = n637 ^ n636 ;
  assign n652 = n635 ^ n619 ;
  assign n653 = n633 ^ n621 ;
  assign n654 = n631 ^ n623 ;
  assign n655 = n611 ^ n607 ;
  assign n656 = n606 ^ n602 ;
  assign n657 = n593 ^ n592 ;
  assign n658 = n595 ^ n594 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = n601 ^ n597 ;
  assign n661 = n659 & n660 ;
  assign n662 = ~n656 & n661 ;
  assign n663 = ~n655 & n662 ;
  assign n664 = n625 ^ x7 ;
  assign n665 = n664 ^ x6 ;
  assign n666 = ~n663 & ~n665 ;
  assign n667 = n626 ^ n624 ;
  assign n668 = n666 & n667 ;
  assign n669 = n627 ^ n559 ;
  assign n670 = ~n668 & n669 ;
  assign n671 = ~n654 & n670 ;
  assign n672 = n632 ^ n622 ;
  assign n673 = ~n671 & ~n672 ;
  assign n674 = n653 & ~n673 ;
  assign n675 = n652 & ~n674 ;
  assign n676 = n651 & ~n675 ;
  assign n638 = ~n636 & ~n637 ;
  assign n618 = n567 ^ n552 ;
  assign n677 = n638 ^ n618 ;
  assign n678 = ~n676 & n677 ;
  assign n617 = n568 ^ n551 ;
  assign n639 = n618 & ~n638 ;
  assign n640 = ~n617 & n639 ;
  assign n616 = n570 ^ n569 ;
  assign n650 = n640 ^ n616 ;
  assign n786 = n678 ^ n650 ;
  assign n691 = n677 ^ n676 ;
  assign n693 = ~x53 & n691 ;
  assign n692 = n691 ^ x53 ;
  assign n694 = n693 ^ n692 ;
  assign n695 = n678 ^ x52 ;
  assign n696 = n675 ^ n651 ;
  assign n697 = n696 ^ x54 ;
  assign n698 = n674 ^ x40 ;
  assign n699 = n669 ^ n668 ;
  assign n700 = n699 ^ x45 ;
  assign n701 = n663 ^ x32 ;
  assign n703 = n658 ^ n657 ;
  assign n704 = n703 ^ x37 ;
  assign n705 = x39 & n592 ;
  assign n706 = n705 ^ n657 ;
  assign n707 = n705 ^ x38 ;
  assign n708 = ~n706 & ~n707 ;
  assign n709 = n708 ^ n658 ;
  assign n710 = ~n704 & ~n709 ;
  assign n702 = n659 ^ x37 ;
  assign n711 = n710 ^ n702 ;
  assign n712 = n659 ^ x36 ;
  assign n713 = n711 & n712 ;
  assign n714 = n713 ^ n660 ;
  assign n717 = n660 ^ n659 ;
  assign n715 = n661 ^ n656 ;
  assign n716 = n715 ^ x35 ;
  assign n718 = n717 ^ n716 ;
  assign n719 = n718 ^ n715 ;
  assign n720 = n714 & ~n719 ;
  assign n721 = n720 ^ n716 ;
  assign n722 = n662 ^ n655 ;
  assign n724 = n722 ^ x34 ;
  assign n723 = n722 ^ n715 ;
  assign n725 = n724 ^ n723 ;
  assign n726 = ~n721 & n725 ;
  assign n727 = n726 ^ n724 ;
  assign n729 = n663 ^ x33 ;
  assign n728 = n722 ^ n663 ;
  assign n730 = n729 ^ n728 ;
  assign n731 = ~n727 & n730 ;
  assign n732 = n731 ^ n729 ;
  assign n733 = n701 & n732 ;
  assign n734 = n733 ^ n665 ;
  assign n737 = n665 ^ n663 ;
  assign n735 = n667 ^ n666 ;
  assign n736 = n735 ^ x47 ;
  assign n738 = n737 ^ n736 ;
  assign n739 = n738 ^ n735 ;
  assign n740 = ~n734 & n739 ;
  assign n741 = n740 ^ n736 ;
  assign n743 = n699 ^ x46 ;
  assign n742 = n735 ^ n699 ;
  assign n744 = n743 ^ n742 ;
  assign n745 = ~n741 & n744 ;
  assign n746 = n745 ^ n743 ;
  assign n747 = n700 & ~n746 ;
  assign n748 = n747 ^ x45 ;
  assign n749 = n748 ^ n670 ;
  assign n750 = n670 ^ x44 ;
  assign n751 = n749 & n750 ;
  assign n752 = n751 ^ n654 ;
  assign n755 = n670 ^ n654 ;
  assign n753 = n672 ^ n671 ;
  assign n754 = n753 ^ x43 ;
  assign n756 = n755 ^ n754 ;
  assign n757 = n756 ^ n753 ;
  assign n758 = ~n752 & n757 ;
  assign n759 = n758 ^ n754 ;
  assign n760 = n673 ^ n653 ;
  assign n762 = n760 ^ x42 ;
  assign n761 = n760 ^ n753 ;
  assign n763 = n762 ^ n761 ;
  assign n764 = ~n759 & n763 ;
  assign n765 = n764 ^ n762 ;
  assign n767 = n674 ^ x41 ;
  assign n766 = n760 ^ n674 ;
  assign n768 = n767 ^ n766 ;
  assign n769 = ~n765 & n768 ;
  assign n770 = n769 ^ n767 ;
  assign n771 = n698 & n770 ;
  assign n772 = n771 ^ n652 ;
  assign n775 = n696 ^ x55 ;
  assign n773 = n674 ^ n652 ;
  assign n774 = n773 ^ n696 ;
  assign n776 = n775 ^ n774 ;
  assign n777 = n772 & ~n776 ;
  assign n778 = n777 ^ n775 ;
  assign n779 = n697 & ~n778 ;
  assign n780 = n779 ^ x54 ;
  assign n781 = ~n693 & n780 ;
  assign n782 = n781 ^ n678 ;
  assign n783 = ~n695 & ~n782 ;
  assign n784 = n783 ^ n678 ;
  assign n785 = ~n694 & n784 ;
  assign n787 = n786 ^ n785 ;
  assign n849 = n787 ^ x51 ;
  assign n810 = n734 ^ x47 ;
  assign n811 = n721 ^ x34 ;
  assign n812 = n657 ^ x38 ;
  assign n813 = n812 ^ n705 ;
  assign n814 = n709 ^ x37 ;
  assign n815 = n813 & ~n814 ;
  assign n816 = n711 ^ x36 ;
  assign n817 = ~n815 & n816 ;
  assign n818 = n714 ^ x35 ;
  assign n819 = ~n817 & n818 ;
  assign n820 = n811 & ~n819 ;
  assign n821 = n727 ^ x33 ;
  assign n822 = ~n820 & ~n821 ;
  assign n823 = n732 ^ x32 ;
  assign n824 = ~n822 & n823 ;
  assign n825 = ~n810 & ~n824 ;
  assign n826 = n741 ^ x46 ;
  assign n827 = n825 & ~n826 ;
  assign n828 = n746 ^ x45 ;
  assign n829 = n827 & ~n828 ;
  assign n830 = n750 ^ n748 ;
  assign n831 = ~n829 & n830 ;
  assign n832 = n752 ^ x43 ;
  assign n833 = ~n831 & ~n832 ;
  assign n834 = n759 ^ x42 ;
  assign n835 = n833 & ~n834 ;
  assign n836 = n765 ^ x41 ;
  assign n837 = ~n835 & n836 ;
  assign n838 = n770 ^ x40 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = n772 ^ x55 ;
  assign n841 = n839 & n840 ;
  assign n842 = n778 ^ x54 ;
  assign n843 = n841 & ~n842 ;
  assign n844 = n780 ^ n692 ;
  assign n845 = n843 & n844 ;
  assign n846 = ~n694 & ~n781 ;
  assign n847 = n846 ^ n695 ;
  assign n848 = ~n845 & n847 ;
  assign n866 = n849 ^ n848 ;
  assign n867 = n592 & ~n866 ;
  assign n940 = n867 ^ n866 ;
  assign n941 = x71 & n940 ;
  assign n679 = n650 & ~n678 ;
  assign n641 = ~n616 & ~n640 ;
  assign n648 = n641 ^ n550 ;
  assign n649 = n648 ^ n571 ;
  assign n689 = n679 ^ n649 ;
  assign n789 = n689 ^ x51 ;
  assign n788 = n786 ^ n689 ;
  assign n790 = n789 ^ n788 ;
  assign n791 = n787 & n790 ;
  assign n792 = n791 ^ n789 ;
  assign n851 = n792 ^ x50 ;
  assign n850 = n848 & ~n849 ;
  assign n869 = n851 ^ n850 ;
  assign n868 = n867 ^ n657 ;
  assign n917 = n869 ^ n868 ;
  assign n918 = ~n657 & ~n917 ;
  assign n942 = n941 ^ n918 ;
  assign n943 = n918 ^ x70 ;
  assign n944 = ~n942 & ~n943 ;
  assign n870 = n869 ^ n867 ;
  assign n871 = ~n868 & ~n870 ;
  assign n872 = n871 ^ n657 ;
  assign n919 = n872 ^ n658 ;
  assign n690 = n689 ^ x50 ;
  assign n793 = n690 & ~n792 ;
  assign n794 = n793 ^ x50 ;
  assign n680 = ~n649 & n679 ;
  assign n643 = n572 ^ n549 ;
  assign n642 = n550 & n641 ;
  assign n647 = n643 ^ n642 ;
  assign n684 = n680 ^ n647 ;
  assign n685 = n684 ^ x49 ;
  assign n853 = n794 ^ n685 ;
  assign n852 = n850 & n851 ;
  assign n864 = n853 ^ n852 ;
  assign n920 = n919 ^ n864 ;
  assign n921 = ~n658 & n920 ;
  assign n945 = n944 ^ n921 ;
  assign n878 = n596 ^ n591 ;
  assign n865 = n864 ^ n658 ;
  assign n873 = n872 ^ n864 ;
  assign n874 = ~n865 & n873 ;
  assign n875 = n874 ^ n658 ;
  assign n879 = n878 ^ n875 ;
  assign n686 = ~x49 & n684 ;
  assign n687 = n686 ^ n685 ;
  assign n795 = ~n686 & n794 ;
  assign n855 = ~n687 & ~n795 ;
  assign n681 = n647 & ~n680 ;
  assign n688 = n681 ^ x48 ;
  assign n856 = n855 ^ n688 ;
  assign n854 = ~n852 & n853 ;
  assign n876 = n856 ^ n854 ;
  assign n923 = n879 ^ n876 ;
  assign n924 = ~n878 & ~n923 ;
  assign n922 = ~n918 & ~n921 ;
  assign n938 = n924 ^ n922 ;
  assign n948 = n938 ^ x69 ;
  assign n946 = n921 ^ n918 ;
  assign n947 = n946 ^ n938 ;
  assign n949 = n948 ^ n947 ;
  assign n950 = ~n945 & ~n949 ;
  assign n951 = n950 ^ n948 ;
  assign n1155 = n951 ^ x68 ;
  assign n1150 = n940 ^ x71 ;
  assign n1151 = n942 ^ x70 ;
  assign n1152 = ~n1150 & n1151 ;
  assign n1153 = n945 ^ x69 ;
  assign n1154 = ~n1152 & n1153 ;
  assign n1996 = n1155 ^ n1154 ;
  assign n1227 = n821 ^ n820 ;
  assign n1189 = n818 ^ n817 ;
  assign n1208 = n1189 ^ n651 ;
  assign n1190 = n1189 ^ n652 ;
  assign n1096 = n592 ^ x39 ;
  assign n803 = n575 ^ n546 ;
  assign n614 = n574 ^ n547 ;
  assign n615 = n573 ^ n548 ;
  assign n644 = ~n642 & n643 ;
  assign n645 = n615 & n644 ;
  assign n804 = n614 & n645 ;
  assign n892 = n803 & n804 ;
  assign n891 = n576 ^ n545 ;
  assign n893 = n892 ^ n891 ;
  assign n805 = n804 ^ n803 ;
  assign n646 = n645 ^ n614 ;
  assign n806 = ~n646 & n681 ;
  assign n894 = ~n805 & n806 ;
  assign n902 = ~n893 & n894 ;
  assign n999 = n577 ^ n544 ;
  assign n1000 = n891 & n892 ;
  assign n1001 = n999 & n1000 ;
  assign n998 = n578 ^ n543 ;
  assign n1002 = n1001 ^ n998 ;
  assign n1020 = ~n902 & n1002 ;
  assign n1022 = n579 ^ n542 ;
  assign n1021 = ~n998 & ~n1001 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1050 = ~n1020 & ~n1023 ;
  assign n1048 = n580 ^ n541 ;
  assign n1047 = ~n1021 & ~n1022 ;
  assign n1049 = n1048 ^ n1047 ;
  assign n1051 = n1050 ^ n1049 ;
  assign n1003 = n1002 ^ n902 ;
  assign n975 = ~x60 & n902 ;
  assign n903 = n902 ^ x60 ;
  assign n976 = n975 ^ n903 ;
  assign n895 = n894 ^ n893 ;
  assign n896 = n895 ^ x61 ;
  assign n993 = n895 ^ x62 ;
  assign n807 = n806 ^ n805 ;
  assign n808 = n807 ^ x62 ;
  assign n682 = n681 ^ n646 ;
  assign n683 = n682 ^ x63 ;
  assign n796 = n795 ^ n681 ;
  assign n797 = ~n688 & ~n796 ;
  assign n798 = n797 ^ n681 ;
  assign n799 = ~n687 & n798 ;
  assign n977 = n975 ^ n682 ;
  assign n978 = n977 ^ x63 ;
  assign n979 = ~n799 & ~n978 ;
  assign n988 = n683 & ~n979 ;
  assign n989 = n682 & n988 ;
  assign n990 = n989 ^ n682 ;
  assign n980 = n979 ^ n807 ;
  assign n981 = n980 ^ n683 ;
  assign n982 = n981 ^ n682 ;
  assign n991 = n990 ^ n982 ;
  assign n992 = ~n808 & n991 ;
  assign n994 = n993 ^ n992 ;
  assign n995 = ~n896 & n994 ;
  assign n996 = n995 ^ x61 ;
  assign n997 = ~n976 & ~n996 ;
  assign n1004 = n1003 ^ n997 ;
  assign n1024 = n1023 ^ n1020 ;
  assign n1025 = n1024 ^ x59 ;
  assign n1026 = n1025 ^ n1003 ;
  assign n1027 = n1026 ^ n1024 ;
  assign n1028 = n1004 & n1027 ;
  assign n1029 = n1028 ^ n1025 ;
  assign n1053 = n1051 ^ x58 ;
  assign n1052 = n1051 ^ n1024 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n1055 = ~n1029 & n1054 ;
  assign n1056 = n1055 ^ n1053 ;
  assign n1077 = n1056 ^ n1049 ;
  assign n1078 = n1051 & ~n1077 ;
  assign n1076 = x57 ^ x56 ;
  assign n1079 = n1078 ^ n1076 ;
  assign n1030 = n1029 ^ x58 ;
  assign n1005 = n1004 ^ x59 ;
  assign n800 = n799 ^ n682 ;
  assign n801 = ~n683 & ~n800 ;
  assign n802 = n801 ^ x63 ;
  assign n888 = n807 ^ n802 ;
  assign n889 = ~n808 & n888 ;
  assign n890 = n889 ^ x62 ;
  assign n901 = n895 ^ n890 ;
  assign n906 = n890 ^ x61 ;
  assign n907 = n901 & n906 ;
  assign n904 = n903 ^ x61 ;
  assign n908 = n907 ^ n904 ;
  assign n897 = n896 ^ n890 ;
  assign n809 = n808 ^ n802 ;
  assign n857 = n854 & ~n856 ;
  assign n858 = n799 ^ n683 ;
  assign n859 = ~n857 & n858 ;
  assign n898 = ~n809 & n859 ;
  assign n909 = ~n897 & n898 ;
  assign n1006 = n908 & ~n909 ;
  assign n1031 = ~n1005 & ~n1006 ;
  assign n1058 = ~n1030 & ~n1031 ;
  assign n1073 = n1058 ^ x57 ;
  assign n1074 = n1058 ^ n1056 ;
  assign n1075 = ~n1073 & n1074 ;
  assign n1080 = n1079 ^ n1075 ;
  assign n1097 = n1096 ^ n1080 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1042 = n1032 ^ n667 ;
  assign n899 = n898 ^ n897 ;
  assign n860 = n859 ^ n809 ;
  assign n861 = n860 ^ n656 ;
  assign n862 = n858 ^ n857 ;
  assign n863 = n862 ^ n660 ;
  assign n881 = n876 ^ n862 ;
  assign n877 = n876 ^ n875 ;
  assign n880 = ~n877 & n879 ;
  assign n882 = n881 ^ n880 ;
  assign n883 = ~n863 & n882 ;
  assign n884 = n883 ^ n660 ;
  assign n885 = n884 ^ n860 ;
  assign n886 = n861 & n885 ;
  assign n887 = n886 ^ n656 ;
  assign n900 = n899 ^ n887 ;
  assign n932 = n887 ^ n655 ;
  assign n914 = ~n900 & n932 ;
  assign n910 = n909 ^ n908 ;
  assign n911 = n910 ^ n655 ;
  assign n915 = n914 ^ n911 ;
  assign n613 = n612 ^ x7 ;
  assign n1009 = n910 ^ n613 ;
  assign n1010 = ~n915 & n1009 ;
  assign n1007 = n1006 ^ n1005 ;
  assign n1008 = n1007 ^ n910 ;
  assign n1011 = n1010 ^ n1008 ;
  assign n1016 = n1007 ^ n665 ;
  assign n1017 = ~n1011 & ~n1016 ;
  assign n1018 = n1017 ^ n665 ;
  assign n1043 = n1032 ^ n1018 ;
  assign n1044 = ~n1042 & ~n1043 ;
  assign n1045 = n1044 ^ n667 ;
  assign n1046 = n1045 ^ n669 ;
  assign n1057 = n1056 ^ x57 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1072 = n1059 ^ n1045 ;
  assign n1084 = n1046 & n1072 ;
  assign n1081 = n1080 ^ n669 ;
  assign n1085 = n1084 ^ n1081 ;
  assign n1069 = n630 ^ n561 ;
  assign n1094 = n1080 ^ n1069 ;
  assign n1095 = ~n1085 & n1094 ;
  assign n1098 = n1097 ^ n1095 ;
  assign n1107 = n1096 ^ n654 ;
  assign n1108 = ~n1098 & ~n1107 ;
  assign n1109 = n1108 ^ n1096 ;
  assign n1119 = n1109 ^ n672 ;
  assign n1122 = n1109 ^ n813 ;
  assign n1123 = n1119 & n1122 ;
  assign n1120 = n813 ^ n653 ;
  assign n1124 = n1123 ^ n1120 ;
  assign n1125 = n814 ^ n813 ;
  assign n1138 = n1125 ^ n653 ;
  assign n1139 = ~n1124 & n1138 ;
  assign n1136 = n816 ^ n815 ;
  assign n1137 = n1136 ^ n1125 ;
  assign n1140 = n1139 ^ n1137 ;
  assign n1135 = n634 ^ n620 ;
  assign n1186 = n1136 ^ n1135 ;
  assign n1187 = ~n1140 & n1186 ;
  assign n1188 = n1187 ^ n1136 ;
  assign n1206 = n1188 ^ n652 ;
  assign n1207 = n1190 & n1206 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1210 = n819 ^ n811 ;
  assign n1224 = n1210 ^ n651 ;
  assign n1225 = ~n1209 & ~n1224 ;
  assign n1226 = n1225 ^ n1210 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1913 = n1228 ^ n677 ;
  assign n1211 = n1210 ^ n1209 ;
  assign n1914 = n1913 ^ n1211 ;
  assign n1191 = n1190 ^ n1188 ;
  assign n1870 = n1191 ^ n1150 ;
  assign n1282 = n1226 ^ n677 ;
  assign n1283 = ~n1228 & ~n1282 ;
  assign n1279 = n639 ^ n617 ;
  assign n1280 = n1279 ^ n677 ;
  assign n1284 = n1283 ^ n1280 ;
  assign n1285 = n823 ^ n822 ;
  assign n1311 = n1285 ^ n1279 ;
  assign n1312 = n1284 & ~n1311 ;
  assign n1310 = n1279 ^ n650 ;
  assign n1313 = n1312 ^ n1310 ;
  assign n1314 = n824 ^ n810 ;
  assign n1343 = n1314 ^ n650 ;
  assign n1344 = n1313 & ~n1343 ;
  assign n1345 = n1344 ^ n650 ;
  assign n1381 = n1345 ^ n649 ;
  assign n1347 = n826 ^ n825 ;
  assign n1348 = n1381 ^ n1347 ;
  assign n1349 = ~n649 & ~n1348 ;
  assign n1315 = n1314 ^ n1313 ;
  assign n1316 = n650 & ~n1315 ;
  assign n1286 = n1285 ^ n1284 ;
  assign n1287 = ~n1279 & ~n1286 ;
  assign n1229 = ~n677 & n1228 ;
  assign n1212 = n651 & ~n1211 ;
  assign n1192 = ~n652 & ~n1191 ;
  assign n1141 = n1135 & ~n1140 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1127 = n653 & n1126 ;
  assign n1111 = n672 & n1122 ;
  assign n1099 = ~n654 & n1098 ;
  assign n1086 = n1069 & ~n1085 ;
  assign n1060 = n1059 ^ n1046 ;
  assign n1061 = n669 & ~n1060 ;
  assign n1019 = n1018 ^ n667 ;
  assign n1033 = n1032 ^ n1019 ;
  assign n1034 = ~n667 & n1033 ;
  assign n1012 = n665 & n1011 ;
  assign n916 = ~n613 & ~n915 ;
  assign n925 = n922 & n924 ;
  assign n926 = n660 & n882 ;
  assign n927 = n925 & ~n926 ;
  assign n928 = n884 ^ n656 ;
  assign n929 = n928 ^ n860 ;
  assign n930 = ~n656 & n929 ;
  assign n931 = n927 & ~n930 ;
  assign n933 = n932 ^ n899 ;
  assign n934 = ~n655 & ~n933 ;
  assign n935 = n931 & ~n934 ;
  assign n1013 = n916 & n935 ;
  assign n1035 = ~n1012 & ~n1013 ;
  assign n1062 = ~n1034 & n1035 ;
  assign n1087 = ~n1061 & ~n1062 ;
  assign n1100 = n1086 & n1087 ;
  assign n1112 = ~n1099 & n1100 ;
  assign n1128 = ~n1111 & ~n1112 ;
  assign n1142 = ~n1127 & ~n1128 ;
  assign n1193 = n1141 & n1142 ;
  assign n1213 = ~n1192 & ~n1193 ;
  assign n1230 = ~n1212 & ~n1213 ;
  assign n1288 = ~n1229 & ~n1230 ;
  assign n1317 = n1287 & ~n1288 ;
  assign n1350 = ~n1316 & n1317 ;
  assign n1376 = ~n1349 & n1350 ;
  assign n1377 = n1347 ^ n1345 ;
  assign n1382 = ~n1377 & ~n1381 ;
  assign n1378 = n828 ^ n827 ;
  assign n1379 = n1378 ^ n649 ;
  assign n1383 = n1382 ^ n1379 ;
  assign n1384 = ~n647 & ~n1383 ;
  assign n1422 = ~n1376 & ~n1384 ;
  assign n1414 = n644 ^ n615 ;
  assign n1415 = n830 ^ n829 ;
  assign n1417 = n1415 ^ n647 ;
  assign n1416 = n1415 ^ n1378 ;
  assign n1418 = n1417 ^ n1416 ;
  assign n1419 = n1383 & n1418 ;
  assign n1420 = n1419 ^ n1417 ;
  assign n1421 = n1414 & ~n1420 ;
  assign n1423 = n1422 ^ n1421 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n936 = n935 ^ n916 ;
  assign n937 = n936 ^ x64 ;
  assign n954 = n926 ^ n925 ;
  assign n939 = n938 ^ x68 ;
  assign n952 = ~n939 & n951 ;
  assign n953 = n952 ^ x68 ;
  assign n955 = n954 ^ n953 ;
  assign n1157 = n953 ^ x67 ;
  assign n960 = ~n955 & n1157 ;
  assign n956 = n930 ^ n927 ;
  assign n957 = n956 ^ x67 ;
  assign n961 = n960 ^ n957 ;
  assign n962 = n934 ^ n931 ;
  assign n964 = n962 ^ x66 ;
  assign n963 = n962 ^ n956 ;
  assign n965 = n964 ^ n963 ;
  assign n966 = ~n961 & n965 ;
  assign n967 = n966 ^ n964 ;
  assign n969 = n936 ^ x65 ;
  assign n968 = n962 ^ n936 ;
  assign n970 = n969 ^ n968 ;
  assign n971 = ~n967 & n970 ;
  assign n972 = n971 ^ n969 ;
  assign n973 = ~n937 & n972 ;
  assign n974 = n973 ^ x64 ;
  assign n1015 = n1014 ^ n974 ;
  assign n1166 = n974 ^ x79 ;
  assign n1040 = ~n1015 & n1166 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1037 = n1036 ^ x79 ;
  assign n1041 = n1040 ^ n1037 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1065 = n1063 ^ x78 ;
  assign n1064 = n1063 ^ n1036 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1067 = n1041 & ~n1066 ;
  assign n1068 = n1067 ^ n1065 ;
  assign n1088 = n1087 ^ n1086 ;
  assign n1090 = n1088 ^ x77 ;
  assign n1089 = n1088 ^ n1063 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1092 = n1068 & ~n1091 ;
  assign n1093 = n1092 ^ n1090 ;
  assign n1101 = n1100 ^ n1099 ;
  assign n1103 = n1101 ^ x76 ;
  assign n1102 = n1101 ^ n1088 ;
  assign n1104 = n1103 ^ n1102 ;
  assign n1105 = n1093 & ~n1104 ;
  assign n1106 = n1105 ^ n1103 ;
  assign n1113 = n1112 ^ n1111 ;
  assign n1115 = n1113 ^ x75 ;
  assign n1114 = n1113 ^ n1101 ;
  assign n1116 = n1115 ^ n1114 ;
  assign n1117 = ~n1106 & n1116 ;
  assign n1118 = n1117 ^ n1115 ;
  assign n1129 = n1128 ^ n1127 ;
  assign n1131 = n1129 ^ x74 ;
  assign n1130 = n1129 ^ n1113 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1133 = ~n1118 & n1132 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1143 = n1142 ^ n1141 ;
  assign n1145 = n1143 ^ x73 ;
  assign n1144 = n1143 ^ n1129 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1147 = n1134 & ~n1146 ;
  assign n1148 = n1147 ^ n1145 ;
  assign n1196 = n1143 ^ x72 ;
  assign n1197 = n1148 & ~n1196 ;
  assign n1198 = n1197 ^ x72 ;
  assign n1194 = n1193 ^ n1192 ;
  assign n1205 = n1198 ^ n1194 ;
  assign n1214 = n1213 ^ n1212 ;
  assign n1215 = n1214 ^ x87 ;
  assign n1216 = n1215 ^ n1198 ;
  assign n1217 = n1216 ^ n1214 ;
  assign n1218 = ~n1205 & n1217 ;
  assign n1219 = n1218 ^ n1215 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1233 = n1231 ^ x86 ;
  assign n1232 = n1231 ^ n1214 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1235 = n1219 & ~n1234 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1289 = n1288 ^ n1287 ;
  assign n1291 = n1289 ^ x85 ;
  assign n1290 = n1289 ^ n1231 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1293 = ~n1236 & n1292 ;
  assign n1294 = n1293 ^ n1291 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1320 = n1318 ^ x84 ;
  assign n1319 = n1318 ^ n1289 ;
  assign n1321 = n1320 ^ n1319 ;
  assign n1322 = ~n1294 & n1321 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1351 = n1350 ^ n1349 ;
  assign n1353 = n1351 ^ x83 ;
  assign n1352 = n1351 ^ n1318 ;
  assign n1354 = n1353 ^ n1352 ;
  assign n1355 = ~n1323 & n1354 ;
  assign n1356 = n1355 ^ n1353 ;
  assign n1385 = n1384 ^ n1376 ;
  assign n1387 = n1385 ^ x82 ;
  assign n1386 = n1385 ^ n1351 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1389 = ~n1356 & n1388 ;
  assign n1390 = n1389 ^ n1387 ;
  assign n1410 = n1385 ^ x81 ;
  assign n1411 = ~n1390 & n1410 ;
  assign n1412 = n1411 ^ x81 ;
  assign n1442 = n1423 ^ n1412 ;
  assign n1450 = n1421 & ~n1422 ;
  assign n1476 = n834 ^ n833 ;
  assign n1477 = n1476 ^ n646 ;
  assign n1443 = n1415 ^ n1414 ;
  assign n1444 = n1420 & n1443 ;
  assign n1445 = n1444 ^ n1414 ;
  assign n1478 = n1477 ^ n1445 ;
  assign n1479 = n1478 ^ n1476 ;
  assign n1447 = n832 ^ n831 ;
  assign n1448 = n1479 ^ n1447 ;
  assign n1449 = n646 & ~n1448 ;
  assign n1451 = n1450 ^ n1449 ;
  assign n1452 = n1451 ^ x80 ;
  assign n1453 = n1452 ^ n1412 ;
  assign n1454 = n1453 ^ n1451 ;
  assign n1455 = ~n1442 & n1454 ;
  assign n1456 = n1455 ^ n1452 ;
  assign n1483 = ~n1449 & ~n1450 ;
  assign n1475 = n1447 ^ n1445 ;
  assign n1480 = ~n1475 & n1479 ;
  assign n1481 = n1480 ^ n1477 ;
  assign n1482 = n805 & ~n1481 ;
  assign n1484 = n1483 ^ n1482 ;
  assign n1486 = n1484 ^ x95 ;
  assign n1485 = n1484 ^ n1451 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1488 = ~n1456 & n1487 ;
  assign n1489 = n1488 ^ n1486 ;
  assign n1546 = ~n1482 & n1483 ;
  assign n1539 = n836 ^ n835 ;
  assign n1541 = n1539 ^ n805 ;
  assign n1540 = n1539 ^ n1476 ;
  assign n1542 = n1541 ^ n1540 ;
  assign n1543 = n1481 & ~n1542 ;
  assign n1544 = n1543 ^ n1541 ;
  assign n1545 = n893 & n1544 ;
  assign n1547 = n1546 ^ n1545 ;
  assign n1549 = n1547 ^ x94 ;
  assign n1548 = n1547 ^ n1484 ;
  assign n1550 = n1549 ^ n1548 ;
  assign n1551 = n1489 & ~n1550 ;
  assign n1552 = n1551 ^ n1549 ;
  assign n1596 = ~n1545 & n1546 ;
  assign n1588 = n1000 ^ n999 ;
  assign n1589 = n838 ^ n837 ;
  assign n1591 = n1589 ^ n893 ;
  assign n1590 = n1589 ^ n1539 ;
  assign n1592 = n1591 ^ n1590 ;
  assign n1593 = ~n1544 & n1592 ;
  assign n1594 = n1593 ^ n1591 ;
  assign n1595 = n1588 & n1594 ;
  assign n1597 = n1596 ^ n1595 ;
  assign n1599 = n1597 ^ x93 ;
  assign n1598 = n1597 ^ n1547 ;
  assign n1600 = n1599 ^ n1598 ;
  assign n1601 = n1552 & ~n1600 ;
  assign n1602 = n1601 ^ n1599 ;
  assign n1653 = n1595 & ~n1596 ;
  assign n1704 = n842 ^ n841 ;
  assign n1705 = n1704 ^ n1002 ;
  assign n1646 = n1589 ^ n1588 ;
  assign n1647 = ~n1594 & n1646 ;
  assign n1648 = n1647 ^ n1588 ;
  assign n1706 = n1705 ^ n1648 ;
  assign n1707 = n1706 ^ n1704 ;
  assign n1650 = n840 ^ n839 ;
  assign n1651 = n1707 ^ n1650 ;
  assign n1652 = n1002 & n1651 ;
  assign n1654 = n1653 ^ n1652 ;
  assign n1656 = n1654 ^ x92 ;
  assign n1655 = n1654 ^ n1597 ;
  assign n1657 = n1656 ^ n1655 ;
  assign n1658 = ~n1602 & n1657 ;
  assign n1659 = n1658 ^ n1656 ;
  assign n1711 = ~n1652 & n1653 ;
  assign n1703 = n1650 ^ n1648 ;
  assign n1708 = ~n1703 & ~n1707 ;
  assign n1709 = n1708 ^ n1705 ;
  assign n1710 = n1023 & n1709 ;
  assign n1712 = n1711 ^ n1710 ;
  assign n1714 = n1712 ^ x91 ;
  assign n1713 = n1712 ^ n1654 ;
  assign n1715 = n1714 ^ n1713 ;
  assign n1716 = ~n1659 & n1715 ;
  assign n1717 = n1716 ^ n1714 ;
  assign n1718 = n1717 ^ x90 ;
  assign n1660 = n1659 ^ x91 ;
  assign n1603 = n1602 ^ x92 ;
  assign n1553 = n1552 ^ x93 ;
  assign n1490 = n1489 ^ x94 ;
  assign n1457 = n1456 ^ x95 ;
  assign n1424 = n1454 ^ n1423 ;
  assign n1391 = n1390 ^ x81 ;
  assign n1357 = n1356 ^ x82 ;
  assign n1324 = n1323 ^ x83 ;
  assign n1295 = n1294 ^ x84 ;
  assign n1237 = n1236 ^ x85 ;
  assign n1220 = n1219 ^ x86 ;
  assign n1195 = n1194 ^ x87 ;
  assign n1199 = n1198 ^ n1195 ;
  assign n1149 = n1148 ^ x72 ;
  assign n1156 = ~n1154 & n1155 ;
  assign n1158 = n1157 ^ n954 ;
  assign n1159 = n1156 & ~n1158 ;
  assign n1160 = n961 ^ x66 ;
  assign n1161 = ~n1159 & n1160 ;
  assign n1162 = n967 ^ x65 ;
  assign n1163 = ~n1161 & ~n1162 ;
  assign n1164 = n972 ^ x64 ;
  assign n1165 = n1163 & n1164 ;
  assign n1167 = n1166 ^ n1014 ;
  assign n1168 = ~n1165 & n1167 ;
  assign n1169 = n1041 ^ x78 ;
  assign n1170 = n1168 & ~n1169 ;
  assign n1171 = n1068 ^ x77 ;
  assign n1172 = n1170 & ~n1171 ;
  assign n1173 = n1093 ^ x76 ;
  assign n1174 = n1172 & ~n1173 ;
  assign n1175 = n1106 ^ x75 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1177 = n1118 ^ x74 ;
  assign n1178 = n1176 & ~n1177 ;
  assign n1179 = n1134 ^ x73 ;
  assign n1180 = n1178 & n1179 ;
  assign n1200 = ~n1149 & ~n1180 ;
  assign n1221 = n1199 & n1200 ;
  assign n1238 = ~n1220 & n1221 ;
  assign n1296 = n1237 & n1238 ;
  assign n1325 = n1295 & n1296 ;
  assign n1358 = n1324 & n1325 ;
  assign n1392 = ~n1357 & ~n1358 ;
  assign n1425 = n1391 & ~n1392 ;
  assign n1458 = n1424 & n1425 ;
  assign n1491 = n1457 & n1458 ;
  assign n1554 = ~n1490 & n1491 ;
  assign n1604 = n1553 & ~n1554 ;
  assign n1661 = n1603 & ~n1604 ;
  assign n1719 = n1660 & n1661 ;
  assign n1765 = ~n1718 & ~n1719 ;
  assign n1773 = ~n1710 & ~n1711 ;
  assign n1766 = n844 ^ n843 ;
  assign n1768 = n1766 ^ n1023 ;
  assign n1767 = n1766 ^ n1704 ;
  assign n1769 = n1768 ^ n1767 ;
  assign n1770 = ~n1709 & ~n1769 ;
  assign n1771 = n1770 ^ n1768 ;
  assign n1772 = n1049 & n1771 ;
  assign n1774 = n1773 ^ n1772 ;
  assign n1776 = n1774 ^ x90 ;
  assign n1775 = n1774 ^ n1712 ;
  assign n1777 = n1776 ^ n1775 ;
  assign n1778 = ~n1717 & n1777 ;
  assign n1779 = n1778 ^ n1776 ;
  assign n1780 = n1779 ^ x89 ;
  assign n1839 = ~n1765 & ~n1780 ;
  assign n1826 = n1047 ^ n541 ;
  assign n1827 = n1048 & n1826 ;
  assign n1828 = n1827 ^ n581 ;
  assign n1832 = n1766 ^ n1049 ;
  assign n1833 = ~n1771 & n1832 ;
  assign n1829 = n1828 ^ n845 ;
  assign n1830 = n1829 ^ n847 ;
  assign n1831 = n1830 ^ n1049 ;
  assign n1834 = n1833 ^ n1831 ;
  assign n1835 = n1828 & ~n1834 ;
  assign n1825 = x89 ^ x88 ;
  assign n1836 = n1835 ^ n1825 ;
  assign n1824 = ~n1772 & n1773 ;
  assign n1837 = n1836 ^ n1824 ;
  assign n1822 = n1774 ^ x89 ;
  assign n1823 = n1779 & ~n1822 ;
  assign n1838 = n1837 ^ n1823 ;
  assign n1840 = n1839 ^ n1838 ;
  assign n1781 = n1780 ^ n1765 ;
  assign n1763 = n1140 ^ n1135 ;
  assign n1817 = n1781 ^ n1763 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1759 = n1720 ^ n1126 ;
  assign n1662 = n1661 ^ n1660 ;
  assign n1644 = n1122 ^ n672 ;
  assign n1698 = n1662 ^ n1644 ;
  assign n1605 = n1604 ^ n1603 ;
  assign n1586 = n1098 ^ n654 ;
  assign n1640 = n1605 ^ n1586 ;
  assign n1555 = n1554 ^ n1553 ;
  assign n1537 = n1085 ^ n1069 ;
  assign n1582 = n1555 ^ n1537 ;
  assign n1492 = n1491 ^ n1490 ;
  assign n1533 = n1492 ^ n1060 ;
  assign n1459 = n1458 ^ n1457 ;
  assign n1470 = n1459 ^ n1033 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n1408 = n1011 ^ n665 ;
  assign n1437 = n1426 ^ n1408 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n1374 = n915 ^ n613 ;
  assign n1404 = n1393 ^ n1374 ;
  assign n1359 = n1358 ^ n1357 ;
  assign n1370 = n1359 ^ n933 ;
  assign n1326 = n1325 ^ n1324 ;
  assign n1297 = n1296 ^ n1295 ;
  assign n1327 = n1326 ^ n1297 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1181 = n1180 ^ n1149 ;
  assign n1182 = n866 ^ n592 ;
  assign n1184 = n1181 & ~n1182 ;
  assign n1185 = n1184 ^ n917 ;
  assign n1201 = n1200 ^ n1199 ;
  assign n1202 = n1201 ^ n1184 ;
  assign n1203 = ~n1185 & ~n1202 ;
  assign n1204 = n1203 ^ n917 ;
  assign n1223 = n1222 ^ n1204 ;
  assign n1255 = n1204 ^ n920 ;
  assign n1243 = ~n1223 & ~n1255 ;
  assign n1239 = n1238 ^ n1237 ;
  assign n1240 = n1239 ^ n920 ;
  assign n1244 = n1243 ^ n1240 ;
  assign n1275 = n1239 ^ n923 ;
  assign n1276 = ~n1244 & ~n1275 ;
  assign n1277 = n1276 ^ n923 ;
  assign n1274 = n882 ^ n660 ;
  assign n1278 = n1277 ^ n1274 ;
  assign n1308 = n1297 ^ n1277 ;
  assign n1309 = ~n1278 & ~n1308 ;
  assign n1328 = n1327 ^ n1309 ;
  assign n1339 = n1326 ^ n929 ;
  assign n1340 = ~n1328 & n1339 ;
  assign n1341 = n1340 ^ n929 ;
  assign n1371 = n1359 ^ n1341 ;
  assign n1372 = n1370 & n1371 ;
  assign n1373 = n1372 ^ n933 ;
  assign n1405 = n1393 ^ n1373 ;
  assign n1406 = n1404 & ~n1405 ;
  assign n1407 = n1406 ^ n1374 ;
  assign n1438 = n1426 ^ n1407 ;
  assign n1439 = ~n1437 & n1438 ;
  assign n1440 = n1439 ^ n1408 ;
  assign n1471 = n1459 ^ n1440 ;
  assign n1472 = n1470 & n1471 ;
  assign n1473 = n1472 ^ n1033 ;
  assign n1534 = n1492 ^ n1473 ;
  assign n1535 = n1533 & n1534 ;
  assign n1536 = n1535 ^ n1060 ;
  assign n1583 = n1555 ^ n1536 ;
  assign n1584 = n1582 & n1583 ;
  assign n1585 = n1584 ^ n1537 ;
  assign n1641 = n1605 ^ n1585 ;
  assign n1642 = ~n1640 & n1641 ;
  assign n1643 = n1642 ^ n1586 ;
  assign n1699 = n1662 ^ n1643 ;
  assign n1700 = ~n1698 & ~n1699 ;
  assign n1701 = n1700 ^ n1644 ;
  assign n1760 = n1720 ^ n1701 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = n1761 ^ n1126 ;
  assign n1818 = n1781 ^ n1762 ;
  assign n1819 = n1817 & ~n1818 ;
  assign n1820 = n1819 ^ n1763 ;
  assign n1867 = n1840 ^ n1820 ;
  assign n1868 = n1840 ^ n1191 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1871 = n1870 ^ n1869 ;
  assign n1911 = n1211 ^ n1150 ;
  assign n1912 = ~n1871 & n1911 ;
  assign n1915 = n1914 ^ n1912 ;
  assign n1910 = n1151 ^ n1150 ;
  assign n1952 = n1913 ^ n1910 ;
  assign n1953 = ~n1915 & n1952 ;
  assign n1950 = n1913 ^ n1286 ;
  assign n1954 = n1953 ^ n1950 ;
  assign n1992 = n1315 ^ n1286 ;
  assign n1955 = n1153 ^ n1152 ;
  assign n1991 = n1955 ^ n1315 ;
  assign n1993 = n1992 ^ n1991 ;
  assign n1994 = ~n1954 & n1993 ;
  assign n1995 = n1994 ^ n1992 ;
  assign n1997 = n1996 ^ n1995 ;
  assign n1998 = n1315 ^ n650 ;
  assign n1999 = n1997 & ~n1998 ;
  assign n2000 = n1999 ^ n650 ;
  assign n1956 = n1955 ^ n1954 ;
  assign n1957 = n1286 ^ n1279 ;
  assign n1958 = n1956 & ~n1957 ;
  assign n1959 = n1958 ^ n1279 ;
  assign n1916 = n1915 ^ n1910 ;
  assign n1917 = n1228 & ~n1916 ;
  assign n1918 = n1917 ^ n677 ;
  assign n1866 = n1211 ^ n651 ;
  assign n1872 = n1871 ^ n1211 ;
  assign n1873 = ~n1866 & ~n1872 ;
  assign n1874 = n1873 ^ n651 ;
  assign n1816 = n1189 ^ n1188 ;
  assign n1821 = n1820 ^ n1191 ;
  assign n1841 = n1840 ^ n1821 ;
  assign n1842 = ~n1816 & ~n1841 ;
  assign n1843 = n1842 ^ n652 ;
  assign n1764 = n1763 ^ n1762 ;
  assign n1782 = n1781 ^ n1764 ;
  assign n1783 = ~n1140 & n1782 ;
  assign n1784 = n1783 ^ n1135 ;
  assign n1697 = n1126 ^ n653 ;
  assign n1702 = n1701 ^ n1126 ;
  assign n1721 = n1720 ^ n1702 ;
  assign n1722 = n1697 & n1721 ;
  assign n1723 = n1722 ^ n653 ;
  assign n1645 = n1644 ^ n1643 ;
  assign n1663 = n1662 ^ n1645 ;
  assign n1664 = n1122 & ~n1663 ;
  assign n1665 = n1664 ^ n672 ;
  assign n1587 = n1586 ^ n1585 ;
  assign n1606 = n1605 ^ n1587 ;
  assign n1607 = ~n1098 & ~n1606 ;
  assign n1608 = n1607 ^ n654 ;
  assign n1538 = n1537 ^ n1536 ;
  assign n1556 = n1555 ^ n1538 ;
  assign n1557 = ~n1085 & ~n1556 ;
  assign n1558 = n1557 ^ n1069 ;
  assign n1474 = n1473 ^ n1060 ;
  assign n1493 = n1492 ^ n1474 ;
  assign n1494 = ~n1072 & n1493 ;
  assign n1495 = n1494 ^ n669 ;
  assign n1441 = n1440 ^ n1033 ;
  assign n1460 = n1459 ^ n1441 ;
  assign n1461 = n1043 & ~n1460 ;
  assign n1462 = n1461 ^ n667 ;
  assign n1409 = n1408 ^ n1407 ;
  assign n1427 = n1426 ^ n1409 ;
  assign n1428 = n1011 & n1427 ;
  assign n1429 = n1428 ^ n665 ;
  assign n1375 = n1374 ^ n1373 ;
  assign n1394 = n1393 ^ n1375 ;
  assign n1395 = ~n915 & ~n1394 ;
  assign n1396 = n1395 ^ n613 ;
  assign n1342 = n1341 ^ n933 ;
  assign n1360 = n1359 ^ n1342 ;
  assign n1361 = n900 & n1360 ;
  assign n1362 = n1361 ^ n655 ;
  assign n1329 = n1328 ^ n929 ;
  assign n1330 = ~n885 & n1329 ;
  assign n1331 = n1330 ^ n656 ;
  assign n1298 = n1297 ^ n1278 ;
  assign n1299 = ~n882 & n1298 ;
  assign n1300 = n1299 ^ n660 ;
  assign n1245 = n1244 ^ n923 ;
  assign n1246 = ~n877 & ~n1245 ;
  assign n1247 = n1246 ^ n878 ;
  assign n1248 = n1181 ^ n592 ;
  assign n1249 = ~n866 & ~n1248 ;
  assign n1250 = n1249 ^ n592 ;
  assign n1251 = n1201 ^ n1185 ;
  assign n1252 = n870 & ~n1251 ;
  assign n1253 = n1252 ^ n657 ;
  assign n1254 = n1250 & ~n1253 ;
  assign n1256 = n1255 ^ n1222 ;
  assign n1257 = ~n873 & n1256 ;
  assign n1258 = n1257 ^ n658 ;
  assign n1259 = n1254 & ~n1258 ;
  assign n1301 = ~n1247 & ~n1259 ;
  assign n1332 = n1300 & ~n1301 ;
  assign n1363 = ~n1331 & n1332 ;
  assign n1397 = ~n1362 & n1363 ;
  assign n1430 = ~n1396 & ~n1397 ;
  assign n1463 = n1429 & n1430 ;
  assign n1496 = ~n1462 & n1463 ;
  assign n1559 = n1495 & ~n1496 ;
  assign n1609 = n1558 & ~n1559 ;
  assign n1666 = ~n1608 & ~n1609 ;
  assign n1724 = n1665 & ~n1666 ;
  assign n1785 = n1723 & ~n1724 ;
  assign n1844 = n1784 & ~n1785 ;
  assign n1875 = ~n1843 & n1844 ;
  assign n1919 = n1874 & ~n1875 ;
  assign n1960 = ~n1918 & ~n1919 ;
  assign n2001 = ~n1959 & n1960 ;
  assign n2036 = n2000 & ~n2001 ;
  assign n2042 = n1158 ^ n1156 ;
  assign n2038 = n1348 ^ n1315 ;
  assign n2037 = n1996 ^ n1348 ;
  assign n2039 = n2038 ^ n2037 ;
  assign n2040 = n1995 & ~n2039 ;
  assign n2041 = n2040 ^ n2038 ;
  assign n2043 = n2042 ^ n2041 ;
  assign n2044 = n1377 & n2043 ;
  assign n2045 = n2044 ^ n649 ;
  assign n2086 = n2036 & ~n2045 ;
  assign n2082 = n1160 ^ n1159 ;
  assign n2076 = n1383 ^ n647 ;
  assign n2078 = n2076 ^ n1348 ;
  assign n2077 = n2076 ^ n2042 ;
  assign n2079 = n2078 ^ n2077 ;
  assign n2080 = n2041 & ~n2079 ;
  assign n2081 = n2080 ^ n2078 ;
  assign n2083 = n2082 ^ n2081 ;
  assign n2084 = ~n1383 & ~n2083 ;
  assign n2085 = n2084 ^ n647 ;
  assign n2087 = n2086 ^ n2085 ;
  assign n2046 = n2045 ^ n2036 ;
  assign n2071 = n2046 ^ x114 ;
  assign n1261 = n1258 ^ n1254 ;
  assign n1262 = n1261 ^ x101 ;
  assign n1264 = x103 & ~n1250 ;
  assign n1263 = n1253 ^ n1250 ;
  assign n1265 = n1264 ^ n1263 ;
  assign n1268 = n1263 ^ x102 ;
  assign n1269 = n1265 & ~n1268 ;
  assign n1266 = n1261 ^ x102 ;
  assign n1270 = n1269 ^ n1266 ;
  assign n1271 = ~n1262 & n1270 ;
  assign n1272 = n1271 ^ x101 ;
  assign n1260 = n1259 ^ n1247 ;
  assign n1273 = n1272 ^ n1260 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1303 = n1302 ^ x100 ;
  assign n1304 = n1303 ^ n1260 ;
  assign n1305 = n1304 ^ n1302 ;
  assign n1306 = n1273 & ~n1305 ;
  assign n1307 = n1306 ^ n1303 ;
  assign n1333 = n1332 ^ n1331 ;
  assign n1335 = n1333 ^ x99 ;
  assign n1334 = n1333 ^ n1302 ;
  assign n1336 = n1335 ^ n1334 ;
  assign n1337 = n1307 & ~n1336 ;
  assign n1338 = n1337 ^ n1335 ;
  assign n1364 = n1363 ^ n1362 ;
  assign n1366 = n1364 ^ x98 ;
  assign n1365 = n1364 ^ n1333 ;
  assign n1367 = n1366 ^ n1365 ;
  assign n1368 = n1338 & ~n1367 ;
  assign n1369 = n1368 ^ n1366 ;
  assign n1398 = n1397 ^ n1396 ;
  assign n1400 = n1398 ^ x97 ;
  assign n1399 = n1398 ^ n1364 ;
  assign n1401 = n1400 ^ n1399 ;
  assign n1402 = n1369 & ~n1401 ;
  assign n1403 = n1402 ^ n1400 ;
  assign n1431 = n1430 ^ n1429 ;
  assign n1433 = n1431 ^ x96 ;
  assign n1432 = n1431 ^ n1398 ;
  assign n1434 = n1433 ^ n1432 ;
  assign n1435 = n1403 & ~n1434 ;
  assign n1436 = n1435 ^ n1433 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1466 = n1464 ^ x111 ;
  assign n1465 = n1464 ^ n1431 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1468 = n1436 & ~n1467 ;
  assign n1469 = n1468 ^ n1466 ;
  assign n1497 = n1496 ^ n1495 ;
  assign n1499 = n1497 ^ x110 ;
  assign n1498 = n1497 ^ n1464 ;
  assign n1500 = n1499 ^ n1498 ;
  assign n1501 = ~n1469 & n1500 ;
  assign n1502 = n1501 ^ n1499 ;
  assign n1560 = n1559 ^ n1558 ;
  assign n1562 = n1560 ^ x109 ;
  assign n1561 = n1560 ^ n1497 ;
  assign n1563 = n1562 ^ n1561 ;
  assign n1564 = n1502 & ~n1563 ;
  assign n1565 = n1564 ^ n1562 ;
  assign n1610 = n1609 ^ n1608 ;
  assign n1612 = n1610 ^ x108 ;
  assign n1611 = n1610 ^ n1560 ;
  assign n1613 = n1612 ^ n1611 ;
  assign n1614 = ~n1565 & n1613 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1667 = n1666 ^ n1665 ;
  assign n1669 = n1667 ^ x107 ;
  assign n1668 = n1667 ^ n1610 ;
  assign n1670 = n1669 ^ n1668 ;
  assign n1671 = ~n1615 & n1670 ;
  assign n1672 = n1671 ^ n1669 ;
  assign n1727 = n1667 ^ x106 ;
  assign n1728 = ~n1672 & n1727 ;
  assign n1729 = n1728 ^ x106 ;
  assign n1725 = n1724 ^ n1723 ;
  assign n1758 = n1729 ^ n1725 ;
  assign n1786 = n1785 ^ n1784 ;
  assign n1787 = n1786 ^ x105 ;
  assign n1788 = n1787 ^ n1786 ;
  assign n1789 = n1788 ^ n1729 ;
  assign n1790 = n1758 & n1789 ;
  assign n1791 = n1790 ^ n1787 ;
  assign n1847 = n1786 ^ x104 ;
  assign n1848 = ~n1791 & n1847 ;
  assign n1849 = n1848 ^ x104 ;
  assign n1845 = n1844 ^ n1843 ;
  assign n1865 = n1849 ^ n1845 ;
  assign n1876 = n1875 ^ n1874 ;
  assign n1877 = n1876 ^ x119 ;
  assign n1878 = n1877 ^ n1849 ;
  assign n1879 = n1878 ^ n1876 ;
  assign n1880 = ~n1865 & n1879 ;
  assign n1881 = n1880 ^ n1877 ;
  assign n1920 = n1919 ^ n1918 ;
  assign n1922 = n1920 ^ x118 ;
  assign n1921 = n1920 ^ n1876 ;
  assign n1923 = n1922 ^ n1921 ;
  assign n1924 = n1881 & ~n1923 ;
  assign n1925 = n1924 ^ n1922 ;
  assign n1961 = n1960 ^ n1959 ;
  assign n1963 = n1961 ^ x117 ;
  assign n1962 = n1961 ^ n1920 ;
  assign n1964 = n1963 ^ n1962 ;
  assign n1965 = n1925 & ~n1964 ;
  assign n1966 = n1965 ^ n1963 ;
  assign n2002 = n2001 ^ n2000 ;
  assign n2004 = n2002 ^ x116 ;
  assign n2003 = n2002 ^ n1961 ;
  assign n2005 = n2004 ^ n2003 ;
  assign n2006 = ~n1966 & n2005 ;
  assign n2007 = n2006 ^ n2004 ;
  assign n2032 = n2002 ^ x115 ;
  assign n2033 = n2007 & ~n2032 ;
  assign n2034 = n2033 ^ x115 ;
  assign n2072 = n2046 ^ n2034 ;
  assign n2073 = ~n2071 & n2072 ;
  assign n2074 = n2073 ^ x114 ;
  assign n2112 = n2087 ^ n2074 ;
  assign n2123 = ~n2085 & ~n2086 ;
  assign n2119 = n1162 ^ n1161 ;
  assign n2113 = n1420 ^ n1414 ;
  assign n2115 = n2113 ^ n2076 ;
  assign n2114 = n2113 ^ n2082 ;
  assign n2116 = n2115 ^ n2114 ;
  assign n2117 = n2081 & n2116 ;
  assign n2118 = n2117 ^ n2115 ;
  assign n2120 = n2119 ^ n2118 ;
  assign n2121 = ~n1420 & n2120 ;
  assign n2122 = n2121 ^ n1414 ;
  assign n2124 = n2123 ^ n2122 ;
  assign n2125 = n2124 ^ x113 ;
  assign n2126 = n2125 ^ n2074 ;
  assign n2127 = n2126 ^ n2124 ;
  assign n2128 = n2112 & n2127 ;
  assign n2129 = n2128 ^ n2125 ;
  assign n2166 = n2122 & n2123 ;
  assign n2160 = n2119 ^ n2113 ;
  assign n2161 = ~n2118 & ~n2160 ;
  assign n2162 = n2161 ^ n2113 ;
  assign n2158 = n1164 ^ n1163 ;
  assign n2159 = n2158 ^ n1448 ;
  assign n2163 = n2162 ^ n2159 ;
  assign n2164 = n1475 & n2163 ;
  assign n2165 = n2164 ^ n646 ;
  assign n2167 = n2166 ^ n2165 ;
  assign n2169 = n2167 ^ x112 ;
  assign n2168 = n2167 ^ n2124 ;
  assign n2170 = n2169 ^ n2168 ;
  assign n2171 = n2129 & ~n2170 ;
  assign n2172 = n2171 ^ n2169 ;
  assign n2173 = n2172 ^ x127 ;
  assign n2130 = n2129 ^ x112 ;
  assign n2075 = n2074 ^ x113 ;
  assign n2088 = n2087 ^ n2075 ;
  assign n2035 = n2034 ^ x114 ;
  assign n2047 = n2046 ^ n2035 ;
  assign n2008 = n2007 ^ x115 ;
  assign n1967 = n1966 ^ x116 ;
  assign n1926 = n1925 ^ x117 ;
  assign n1882 = n1881 ^ x118 ;
  assign n1846 = n1845 ^ x119 ;
  assign n1850 = n1849 ^ n1846 ;
  assign n1792 = n1791 ^ x104 ;
  assign n1726 = n1725 ^ x105 ;
  assign n1730 = n1729 ^ n1726 ;
  assign n1673 = n1672 ^ x106 ;
  assign n1616 = n1615 ^ x107 ;
  assign n1566 = n1565 ^ x108 ;
  assign n1503 = n1502 ^ x109 ;
  assign n1504 = n1264 ^ x102 ;
  assign n1505 = n1504 ^ n1263 ;
  assign n1506 = n1270 ^ x101 ;
  assign n1507 = n1505 & n1506 ;
  assign n1508 = n1272 ^ x100 ;
  assign n1509 = n1508 ^ n1260 ;
  assign n1510 = n1507 & n1509 ;
  assign n1511 = n1307 ^ x99 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = n1338 ^ x98 ;
  assign n1514 = ~n1512 & n1513 ;
  assign n1515 = n1369 ^ x97 ;
  assign n1516 = n1514 & n1515 ;
  assign n1517 = n1403 ^ x96 ;
  assign n1518 = n1516 & n1517 ;
  assign n1519 = n1436 ^ x111 ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = n1469 ^ x110 ;
  assign n1522 = ~n1520 & ~n1521 ;
  assign n1567 = n1503 & n1522 ;
  assign n1617 = ~n1566 & n1567 ;
  assign n1674 = n1616 & ~n1617 ;
  assign n1731 = n1673 & n1674 ;
  assign n1793 = n1730 & ~n1731 ;
  assign n1851 = ~n1792 & n1793 ;
  assign n1883 = ~n1850 & n1851 ;
  assign n1927 = ~n1882 & ~n1883 ;
  assign n1968 = n1926 & ~n1927 ;
  assign n2009 = ~n1967 & n1968 ;
  assign n2048 = n2008 & n2009 ;
  assign n2089 = n2047 & n2048 ;
  assign n2131 = ~n2088 & ~n2089 ;
  assign n2174 = n2130 & ~n2131 ;
  assign n2210 = n2173 & n2174 ;
  assign n2202 = n2165 & n2166 ;
  assign n2197 = n1167 ^ n1165 ;
  assign n2193 = n2162 ^ n2158 ;
  assign n2194 = n2162 ^ n1448 ;
  assign n2195 = n2193 & ~n2194 ;
  assign n2196 = n2195 ^ n1448 ;
  assign n2198 = n2197 ^ n2196 ;
  assign n2199 = n2198 ^ n805 ;
  assign n2200 = ~n1481 & n2199 ;
  assign n2201 = n2200 ^ n805 ;
  assign n2203 = n2202 ^ n2201 ;
  assign n2205 = n2203 ^ x127 ;
  assign n2204 = n2203 ^ n2167 ;
  assign n2206 = n2205 ^ n2204 ;
  assign n2207 = n2172 & ~n2206 ;
  assign n2208 = n2207 ^ n2205 ;
  assign n2209 = n2208 ^ x126 ;
  assign n2211 = n2210 ^ n2209 ;
  assign n2175 = n2174 ^ n2173 ;
  assign n2188 = n2175 ^ n1721 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2153 = n2132 ^ n1663 ;
  assign n2090 = n2089 ^ n2088 ;
  assign n2107 = n2090 ^ n1606 ;
  assign n2049 = n2048 ^ n2047 ;
  assign n2066 = n2049 ^ n1556 ;
  assign n2010 = n2009 ^ n2008 ;
  assign n2027 = n2010 ^ n1493 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n1986 = n1969 ^ n1460 ;
  assign n1928 = n1927 ^ n1926 ;
  assign n1945 = n1928 ^ n1427 ;
  assign n1852 = n1851 ^ n1850 ;
  assign n1794 = n1793 ^ n1792 ;
  assign n1811 = n1794 ^ n1329 ;
  assign n1732 = n1731 ^ n1730 ;
  assign n1753 = n1732 ^ n1298 ;
  assign n1675 = n1674 ^ n1673 ;
  assign n1692 = n1675 ^ n1245 ;
  assign n1618 = n1617 ^ n1616 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1523 = n1522 ^ n1503 ;
  assign n1569 = ~n1183 & ~n1523 ;
  assign n1570 = n1569 ^ n1251 ;
  assign n1568 = n1567 ^ n1566 ;
  assign n1579 = n1569 ^ n1568 ;
  assign n1580 = ~n1570 & ~n1579 ;
  assign n1581 = n1580 ^ n1251 ;
  assign n1619 = n1618 ^ n1581 ;
  assign n1636 = n1581 ^ n1256 ;
  assign n1637 = ~n1619 & ~n1636 ;
  assign n1638 = n1637 ^ n1256 ;
  assign n1693 = n1675 ^ n1638 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = n1694 ^ n1245 ;
  assign n1754 = n1732 ^ n1695 ;
  assign n1755 = n1753 & n1754 ;
  assign n1756 = n1755 ^ n1298 ;
  assign n1812 = n1794 ^ n1756 ;
  assign n1813 = n1811 & ~n1812 ;
  assign n1814 = n1813 ^ n1329 ;
  assign n1864 = n1852 ^ n1814 ;
  assign n1884 = n1883 ^ n1882 ;
  assign n1885 = n1884 ^ n1360 ;
  assign n1886 = n1885 ^ n1884 ;
  assign n1887 = n1886 ^ n1814 ;
  assign n1888 = ~n1864 & n1887 ;
  assign n1889 = n1888 ^ n1885 ;
  assign n1906 = n1884 ^ n1394 ;
  assign n1907 = ~n1889 & ~n1906 ;
  assign n1908 = n1907 ^ n1394 ;
  assign n1946 = n1928 ^ n1908 ;
  assign n1947 = n1945 & n1946 ;
  assign n1948 = n1947 ^ n1427 ;
  assign n1987 = n1969 ^ n1948 ;
  assign n1988 = ~n1986 & ~n1987 ;
  assign n1989 = n1988 ^ n1460 ;
  assign n2028 = n2010 ^ n1989 ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2030 = n2029 ^ n1493 ;
  assign n2067 = n2049 ^ n2030 ;
  assign n2068 = n2066 & n2067 ;
  assign n2069 = n2068 ^ n1556 ;
  assign n2108 = n2090 ^ n2069 ;
  assign n2109 = ~n2107 & n2108 ;
  assign n2110 = n2109 ^ n1606 ;
  assign n2154 = n2132 ^ n2110 ;
  assign n2155 = ~n2153 & n2154 ;
  assign n2156 = n2155 ^ n1663 ;
  assign n2189 = n2175 ^ n2156 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2191 = n2190 ^ n1721 ;
  assign n2229 = n2211 ^ n2191 ;
  assign n1571 = n1570 ^ n1568 ;
  assign n1572 = n1202 & ~n1571 ;
  assign n1573 = n1572 ^ n917 ;
  assign n1524 = n1523 ^ n1182 ;
  assign n1525 = n1181 & ~n1524 ;
  assign n1526 = n1525 ^ n1182 ;
  assign n1531 = n592 & ~n1526 ;
  assign n1532 = n1531 ^ n657 ;
  assign n1574 = n1573 ^ n1532 ;
  assign n1527 = n1526 ^ n592 ;
  assign n1529 = x135 & ~n1527 ;
  assign n1577 = n1574 ^ n1529 ;
  assign n1578 = n1573 ^ n1531 ;
  assign n1620 = n1619 ^ n1256 ;
  assign n1621 = n1223 & n1620 ;
  assign n1622 = n1621 ^ n920 ;
  assign n1623 = n1622 ^ n657 ;
  assign n1624 = n1623 ^ n1573 ;
  assign n1625 = n1624 ^ n1622 ;
  assign n1626 = n1578 & n1625 ;
  assign n1627 = n1626 ^ n1623 ;
  assign n1628 = n1627 ^ n658 ;
  assign n1629 = n1628 ^ x134 ;
  assign n1630 = n1629 ^ n1574 ;
  assign n1631 = n1630 ^ n1628 ;
  assign n1632 = ~n1577 & n1631 ;
  assign n1633 = n1632 ^ n1629 ;
  assign n1639 = n1638 ^ n1245 ;
  assign n1676 = n1675 ^ n1639 ;
  assign n1677 = n1244 & ~n1676 ;
  assign n1678 = n1677 ^ n923 ;
  assign n1680 = n1678 ^ n658 ;
  assign n1679 = n1678 ^ n1622 ;
  assign n1681 = n1680 ^ n1679 ;
  assign n1682 = n1627 & ~n1681 ;
  assign n1683 = n1682 ^ n1680 ;
  assign n1684 = n1683 ^ n878 ;
  assign n1686 = n1684 ^ x133 ;
  assign n1685 = n1684 ^ n1628 ;
  assign n1687 = n1686 ^ n1685 ;
  assign n1688 = ~n1633 & n1687 ;
  assign n1689 = n1688 ^ n1686 ;
  assign n1696 = n1695 ^ n1298 ;
  assign n1733 = n1732 ^ n1696 ;
  assign n1734 = ~n1308 & ~n1733 ;
  assign n1735 = n1734 ^ n1274 ;
  assign n1737 = n1735 ^ n878 ;
  assign n1736 = n1735 ^ n1678 ;
  assign n1738 = n1737 ^ n1736 ;
  assign n1739 = ~n1683 & ~n1738 ;
  assign n1740 = n1739 ^ n1737 ;
  assign n1741 = n1740 ^ n660 ;
  assign n1743 = n1741 ^ x132 ;
  assign n1742 = n1741 ^ n1684 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1745 = ~n1689 & n1744 ;
  assign n1746 = n1745 ^ n1743 ;
  assign n1757 = n1756 ^ n1329 ;
  assign n1795 = n1794 ^ n1757 ;
  assign n1796 = n1328 & n1795 ;
  assign n1797 = n1796 ^ n929 ;
  assign n1749 = n1735 ^ n660 ;
  assign n1750 = n1740 & ~n1749 ;
  assign n1751 = n1750 ^ n660 ;
  assign n1752 = n1751 ^ n656 ;
  assign n1798 = n1797 ^ n1752 ;
  assign n1800 = n1798 ^ x131 ;
  assign n1799 = n1798 ^ n1741 ;
  assign n1801 = n1800 ^ n1799 ;
  assign n1802 = n1746 & ~n1801 ;
  assign n1803 = n1802 ^ n1800 ;
  assign n1815 = n1814 ^ n1360 ;
  assign n1853 = n1852 ^ n1815 ;
  assign n1854 = ~n1371 & n1853 ;
  assign n1806 = n1797 ^ n656 ;
  assign n1807 = n1797 ^ n1751 ;
  assign n1808 = ~n1806 & ~n1807 ;
  assign n1809 = n1808 ^ n656 ;
  assign n1810 = n1809 ^ n933 ;
  assign n1855 = n1854 ^ n1810 ;
  assign n1856 = n1855 ^ n655 ;
  assign n1858 = n1856 ^ x130 ;
  assign n1857 = n1856 ^ n1798 ;
  assign n1859 = n1858 ^ n1857 ;
  assign n1860 = n1803 & ~n1859 ;
  assign n1861 = n1860 ^ n1858 ;
  assign n1890 = n1889 ^ n1374 ;
  assign n1891 = n1405 & n1890 ;
  assign n1892 = n1891 ^ n1374 ;
  assign n1893 = n1892 ^ n655 ;
  assign n1894 = n1893 ^ n1809 ;
  assign n1895 = n1894 ^ n1892 ;
  assign n1896 = ~n1855 & n1895 ;
  assign n1897 = n1896 ^ n1893 ;
  assign n1898 = n1897 ^ n613 ;
  assign n1900 = n1898 ^ x129 ;
  assign n1899 = n1898 ^ n1856 ;
  assign n1901 = n1900 ^ n1899 ;
  assign n1902 = n1861 & ~n1901 ;
  assign n1903 = n1902 ^ n1900 ;
  assign n1909 = n1908 ^ n1427 ;
  assign n1929 = n1928 ^ n1909 ;
  assign n1930 = ~n1438 & ~n1929 ;
  assign n1931 = n1930 ^ n1408 ;
  assign n1933 = n1931 ^ n613 ;
  assign n1932 = n1931 ^ n1892 ;
  assign n1934 = n1933 ^ n1932 ;
  assign n1935 = ~n1897 & ~n1934 ;
  assign n1936 = n1935 ^ n1933 ;
  assign n1937 = n1936 ^ n665 ;
  assign n1939 = n1937 ^ x128 ;
  assign n1938 = n1937 ^ n1898 ;
  assign n1940 = n1939 ^ n1938 ;
  assign n1941 = ~n1903 & n1940 ;
  assign n1942 = n1941 ^ n1939 ;
  assign n1943 = n1942 ^ x143 ;
  assign n1528 = n1527 ^ x135 ;
  assign n1530 = n1529 ^ x134 ;
  assign n1575 = n1574 ^ n1530 ;
  assign n1576 = n1528 & ~n1575 ;
  assign n1634 = n1633 ^ x133 ;
  assign n1635 = n1576 & ~n1634 ;
  assign n1690 = n1689 ^ x132 ;
  assign n1691 = n1635 & ~n1690 ;
  assign n1747 = n1746 ^ x131 ;
  assign n1748 = ~n1691 & ~n1747 ;
  assign n1804 = n1803 ^ x130 ;
  assign n1805 = ~n1748 & n1804 ;
  assign n1862 = n1861 ^ x129 ;
  assign n1863 = ~n1805 & ~n1862 ;
  assign n1904 = n1903 ^ x128 ;
  assign n1905 = ~n1863 & ~n1904 ;
  assign n3007 = n1943 ^ n1905 ;
  assign n2157 = n2156 ^ n1721 ;
  assign n2176 = n2175 ^ n2157 ;
  assign n2111 = n2110 ^ n1663 ;
  assign n2133 = n2132 ^ n2111 ;
  assign n2984 = n2176 ^ n2133 ;
  assign n2853 = n1929 ^ n1528 ;
  assign n2833 = n1889 ^ n1394 ;
  assign n2834 = n2833 ^ n1528 ;
  assign n2399 = n1997 ^ n1315 ;
  assign n2244 = n2201 & n2202 ;
  assign n2233 = n1481 ^ n805 ;
  assign n2234 = n2233 ^ n2196 ;
  assign n2239 = n2198 & n2234 ;
  assign n2235 = n1169 ^ n1168 ;
  assign n2236 = n2235 ^ n2197 ;
  assign n2240 = n2239 ^ n2236 ;
  assign n2241 = n2240 ^ n893 ;
  assign n2242 = n1544 & n2241 ;
  assign n2243 = n2242 ^ n893 ;
  assign n2245 = n2244 ^ n2243 ;
  assign n2247 = n2245 ^ x126 ;
  assign n2246 = n2245 ^ n2203 ;
  assign n2248 = n2247 ^ n2246 ;
  assign n2249 = n2208 & ~n2248 ;
  assign n2250 = n2249 ^ n2247 ;
  assign n2286 = n2243 & n2244 ;
  assign n2282 = n1171 ^ n1170 ;
  assign n2276 = n1594 ^ n1588 ;
  assign n2278 = n2276 ^ n2235 ;
  assign n2275 = n1544 ^ n893 ;
  assign n2277 = n2276 ^ n2275 ;
  assign n2279 = n2278 ^ n2277 ;
  assign n2280 = n2240 & n2279 ;
  assign n2281 = n2280 ^ n2278 ;
  assign n2283 = n2282 ^ n2281 ;
  assign n2284 = n1594 & ~n2283 ;
  assign n2285 = n2284 ^ n1588 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2289 = n2287 ^ x125 ;
  assign n2288 = n2287 ^ n2245 ;
  assign n2290 = n2289 ^ n2288 ;
  assign n2291 = n2250 & ~n2290 ;
  assign n2292 = n2291 ^ n2289 ;
  assign n2293 = n2292 ^ x124 ;
  assign n2251 = n2250 ^ x125 ;
  assign n2252 = ~n2209 & ~n2210 ;
  assign n2294 = ~n2251 & n2252 ;
  assign n2318 = ~n2293 & n2294 ;
  assign n2328 = n2285 & n2286 ;
  assign n2319 = n1173 ^ n1172 ;
  assign n2321 = n2319 ^ n2276 ;
  assign n2320 = n2319 ^ n2282 ;
  assign n2322 = n2321 ^ n2320 ;
  assign n2323 = n2281 & n2322 ;
  assign n2324 = n2323 ^ n2321 ;
  assign n2325 = n2324 ^ n1651 ;
  assign n2326 = n1703 & n2325 ;
  assign n2327 = n2326 ^ n1002 ;
  assign n2329 = n2328 ^ n2327 ;
  assign n2331 = n2329 ^ x124 ;
  assign n2330 = n2329 ^ n2287 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2333 = n2292 & ~n2332 ;
  assign n2334 = n2333 ^ n2331 ;
  assign n2335 = n2334 ^ x123 ;
  assign n2354 = n2318 & ~n2335 ;
  assign n2365 = n2327 & ~n2328 ;
  assign n2361 = n1175 ^ n1174 ;
  assign n2355 = n1709 ^ n1023 ;
  assign n2357 = n2355 ^ n1651 ;
  assign n2356 = n2355 ^ n2319 ;
  assign n2358 = n2357 ^ n2356 ;
  assign n2359 = ~n2324 & ~n2358 ;
  assign n2360 = n2359 ^ n2357 ;
  assign n2362 = n2361 ^ n2360 ;
  assign n2363 = n1709 & n2362 ;
  assign n2364 = n2363 ^ n1023 ;
  assign n2366 = n2365 ^ n2364 ;
  assign n2368 = n2366 ^ x123 ;
  assign n2367 = n2366 ^ n2329 ;
  assign n2369 = n2368 ^ n2367 ;
  assign n2370 = n2334 & ~n2369 ;
  assign n2371 = n2370 ^ n2368 ;
  assign n2372 = n2371 ^ x122 ;
  assign n2422 = n2354 & n2372 ;
  assign n2414 = n2364 & ~n2365 ;
  assign n2410 = n1177 ^ n1176 ;
  assign n2404 = n1771 ^ n1049 ;
  assign n2406 = n2404 ^ n2355 ;
  assign n2405 = n2404 ^ n2361 ;
  assign n2407 = n2406 ^ n2405 ;
  assign n2408 = ~n2360 & n2407 ;
  assign n2409 = n2408 ^ n2406 ;
  assign n2411 = n2410 ^ n2409 ;
  assign n2412 = n1771 & n2411 ;
  assign n2413 = n2412 ^ n1049 ;
  assign n2415 = n2414 ^ n2413 ;
  assign n2417 = n2415 ^ x122 ;
  assign n2416 = n2415 ^ n2366 ;
  assign n2418 = n2417 ^ n2416 ;
  assign n2419 = ~n2371 & n2418 ;
  assign n2420 = n2419 ^ n2417 ;
  assign n2421 = n2420 ^ x121 ;
  assign n2423 = n2422 ^ n2421 ;
  assign n2336 = n2335 ^ n2318 ;
  assign n2374 = n2336 ^ n1916 ;
  assign n2253 = n2252 ^ n2251 ;
  assign n2228 = n2211 ^ n1782 ;
  assign n2230 = n2228 & ~n2229 ;
  assign n2231 = n2230 ^ n1782 ;
  assign n2274 = n2253 ^ n2231 ;
  assign n2295 = n2294 ^ n2293 ;
  assign n2296 = n2295 ^ n1841 ;
  assign n2297 = n2296 ^ n2295 ;
  assign n2298 = n2297 ^ n2231 ;
  assign n2299 = n2274 & ~n2298 ;
  assign n2300 = n2299 ^ n2296 ;
  assign n2314 = n2295 ^ n1872 ;
  assign n2315 = ~n2300 & n2314 ;
  assign n2316 = n2315 ^ n1872 ;
  assign n2375 = n2336 ^ n2316 ;
  assign n2376 = n2374 & ~n2375 ;
  assign n2377 = n2376 ^ n1916 ;
  assign n2378 = n2377 ^ n1956 ;
  assign n2373 = n2372 ^ n2354 ;
  assign n2400 = n2377 ^ n2373 ;
  assign n2401 = ~n2378 & n2400 ;
  assign n2402 = n2401 ^ n1956 ;
  assign n2403 = n2402 ^ n1997 ;
  assign n2424 = n2423 ^ n2403 ;
  assign n2425 = ~n2399 & n2424 ;
  assign n2426 = n2425 ^ n1315 ;
  assign n2301 = n2300 ^ n1211 ;
  assign n2302 = n1871 & n2301 ;
  assign n2303 = n2302 ^ n1211 ;
  assign n2177 = n1760 & n2176 ;
  assign n2178 = n2177 ^ n1126 ;
  assign n1949 = n1948 ^ n1460 ;
  assign n1970 = n1969 ^ n1949 ;
  assign n1971 = ~n1471 & ~n1970 ;
  assign n1972 = n1971 ^ n1033 ;
  assign n1974 = n1972 ^ n665 ;
  assign n1973 = n1972 ^ n1931 ;
  assign n1975 = n1974 ^ n1973 ;
  assign n1976 = n1936 & n1975 ;
  assign n1977 = n1976 ^ n1974 ;
  assign n1990 = n1989 ^ n1493 ;
  assign n2011 = n2010 ^ n1990 ;
  assign n2012 = ~n1534 & n2011 ;
  assign n2013 = n2012 ^ n1060 ;
  assign n2015 = n2013 ^ n667 ;
  assign n2014 = n2013 ^ n1972 ;
  assign n2016 = n2015 ^ n2014 ;
  assign n2017 = n1977 & n2016 ;
  assign n2018 = n2017 ^ n2015 ;
  assign n2031 = n2030 ^ n1556 ;
  assign n2050 = n2049 ^ n2031 ;
  assign n2051 = ~n1583 & n2050 ;
  assign n2052 = n2051 ^ n1537 ;
  assign n2054 = n2052 ^ n669 ;
  assign n2053 = n2052 ^ n2013 ;
  assign n2055 = n2054 ^ n2053 ;
  assign n2056 = n2018 & ~n2055 ;
  assign n2057 = n2056 ^ n2054 ;
  assign n2070 = n2069 ^ n1606 ;
  assign n2091 = n2090 ^ n2070 ;
  assign n2092 = ~n1641 & n2091 ;
  assign n2093 = n2092 ^ n1586 ;
  assign n2095 = n2093 ^ n1069 ;
  assign n2094 = n2093 ^ n2052 ;
  assign n2096 = n2095 ^ n2094 ;
  assign n2097 = ~n2057 & ~n2096 ;
  assign n2098 = n2097 ^ n2095 ;
  assign n2134 = n1699 & n2133 ;
  assign n2135 = n2134 ^ n1644 ;
  assign n2137 = n2135 ^ n654 ;
  assign n2136 = n2135 ^ n2093 ;
  assign n2138 = n2137 ^ n2136 ;
  assign n2139 = n2098 & ~n2138 ;
  assign n2140 = n2139 ^ n2137 ;
  assign n2149 = n2135 ^ n672 ;
  assign n2150 = ~n2140 & n2149 ;
  assign n2151 = n2150 ^ n672 ;
  assign n2187 = n2178 ^ n2151 ;
  assign n2192 = n2191 ^ n1782 ;
  assign n2212 = n2211 ^ n2192 ;
  assign n2213 = n1818 & n2212 ;
  assign n2214 = n2213 ^ n1763 ;
  assign n2215 = n2214 ^ n653 ;
  assign n2216 = n2215 ^ n2151 ;
  assign n2217 = n2216 ^ n2214 ;
  assign n2218 = n2187 & ~n2217 ;
  assign n2219 = n2218 ^ n2215 ;
  assign n2232 = n2231 ^ n1841 ;
  assign n2254 = n2253 ^ n2232 ;
  assign n2255 = n1867 & n2254 ;
  assign n2256 = n2255 ^ n1191 ;
  assign n2258 = n2256 ^ n1135 ;
  assign n2257 = n2256 ^ n2214 ;
  assign n2259 = n2258 ^ n2257 ;
  assign n2260 = ~n2219 & ~n2259 ;
  assign n2261 = n2260 ^ n2258 ;
  assign n2270 = n2256 ^ n652 ;
  assign n2271 = ~n2261 & ~n2270 ;
  assign n2272 = n2271 ^ n652 ;
  assign n2312 = n2303 ^ n2272 ;
  assign n2313 = n1916 ^ n1913 ;
  assign n2317 = n2316 ^ n1916 ;
  assign n2337 = n2336 ^ n2317 ;
  assign n2338 = ~n2313 & ~n2337 ;
  assign n2339 = n2338 ^ n1913 ;
  assign n2340 = n2339 ^ n651 ;
  assign n2341 = n2340 ^ n2303 ;
  assign n2342 = n2341 ^ n2339 ;
  assign n2343 = n2312 & ~n2342 ;
  assign n2344 = n2343 ^ n2340 ;
  assign n2353 = n1956 ^ n1286 ;
  assign n2379 = n2378 ^ n2373 ;
  assign n2380 = ~n2353 & ~n2379 ;
  assign n2381 = n2380 ^ n1286 ;
  assign n2383 = n2381 ^ n677 ;
  assign n2382 = n2381 ^ n2339 ;
  assign n2384 = n2383 ^ n2382 ;
  assign n2385 = ~n2344 & n2384 ;
  assign n2386 = n2385 ^ n2383 ;
  assign n2395 = n2381 ^ n1279 ;
  assign n2396 = n2386 & ~n2395 ;
  assign n2397 = n2396 ^ n1279 ;
  assign n2439 = n2426 ^ n2397 ;
  assign n2440 = n2043 ^ n1348 ;
  assign n2462 = n2421 & ~n2422 ;
  assign n2457 = x121 ^ x120 ;
  assign n2458 = n2457 ^ n1828 ;
  assign n2456 = n2413 & n2414 ;
  assign n2459 = n2458 ^ n2456 ;
  assign n2448 = n1834 ^ n1828 ;
  assign n2452 = n2410 ^ n2404 ;
  assign n2453 = ~n2409 & ~n2452 ;
  assign n2449 = n1834 ^ n1178 ;
  assign n2450 = n2449 ^ n1179 ;
  assign n2451 = n2450 ^ n2410 ;
  assign n2454 = n2453 ^ n2451 ;
  assign n2455 = n2448 & n2454 ;
  assign n2460 = n2459 ^ n2455 ;
  assign n2446 = n2415 ^ x121 ;
  assign n2447 = n2420 & ~n2446 ;
  assign n2461 = n2460 ^ n2447 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2441 = n2423 ^ n1997 ;
  assign n2442 = n2423 ^ n2402 ;
  assign n2443 = n2441 & ~n2442 ;
  assign n2444 = n2443 ^ n1997 ;
  assign n2445 = n2444 ^ n2043 ;
  assign n2464 = n2463 ^ n2445 ;
  assign n2465 = ~n2440 & ~n2464 ;
  assign n2466 = n2465 ^ n1348 ;
  assign n2467 = n2466 ^ n650 ;
  assign n2468 = n2467 ^ n2397 ;
  assign n2469 = n2468 ^ n2466 ;
  assign n2470 = n2439 & n2469 ;
  assign n2471 = n2470 ^ n2467 ;
  assign n2472 = n2471 ^ n649 ;
  assign n1978 = n1977 ^ n667 ;
  assign n1980 = n1978 ^ x143 ;
  assign n1979 = n1978 ^ n1937 ;
  assign n1981 = n1980 ^ n1979 ;
  assign n1982 = ~n1942 & n1981 ;
  assign n1983 = n1982 ^ n1980 ;
  assign n2019 = n2018 ^ n669 ;
  assign n2021 = n2019 ^ x142 ;
  assign n2020 = n2019 ^ n1978 ;
  assign n2022 = n2021 ^ n2020 ;
  assign n2023 = n1983 & ~n2022 ;
  assign n2024 = n2023 ^ n2021 ;
  assign n2058 = n2057 ^ n1069 ;
  assign n2060 = n2058 ^ x141 ;
  assign n2059 = n2058 ^ n2019 ;
  assign n2061 = n2060 ^ n2059 ;
  assign n2062 = n2024 & ~n2061 ;
  assign n2063 = n2062 ^ n2060 ;
  assign n2099 = n2098 ^ n654 ;
  assign n2101 = n2099 ^ x140 ;
  assign n2100 = n2099 ^ n2058 ;
  assign n2102 = n2101 ^ n2100 ;
  assign n2103 = n2063 & ~n2102 ;
  assign n2104 = n2103 ^ n2101 ;
  assign n2141 = n2140 ^ n672 ;
  assign n2143 = n2141 ^ x139 ;
  assign n2142 = n2141 ^ n2099 ;
  assign n2144 = n2143 ^ n2142 ;
  assign n2145 = ~n2104 & n2144 ;
  assign n2146 = n2145 ^ n2143 ;
  assign n2152 = n2151 ^ n653 ;
  assign n2179 = n2178 ^ n2152 ;
  assign n2181 = n2179 ^ x138 ;
  assign n2180 = n2179 ^ n2141 ;
  assign n2182 = n2181 ^ n2180 ;
  assign n2183 = n2146 & ~n2182 ;
  assign n2184 = n2183 ^ n2181 ;
  assign n2220 = n2219 ^ n1135 ;
  assign n2222 = n2220 ^ x137 ;
  assign n2221 = n2220 ^ n2179 ;
  assign n2223 = n2222 ^ n2221 ;
  assign n2224 = n2184 & ~n2223 ;
  assign n2225 = n2224 ^ n2222 ;
  assign n2262 = n2261 ^ n652 ;
  assign n2264 = n2262 ^ x136 ;
  assign n2263 = n2262 ^ n2220 ;
  assign n2265 = n2264 ^ n2263 ;
  assign n2266 = n2225 & ~n2265 ;
  assign n2267 = n2266 ^ n2264 ;
  assign n2273 = n2272 ^ n651 ;
  assign n2304 = n2303 ^ n2273 ;
  assign n2306 = n2304 ^ x151 ;
  assign n2305 = n2304 ^ n2262 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2308 = ~n2267 & n2307 ;
  assign n2309 = n2308 ^ n2306 ;
  assign n2345 = n2344 ^ n677 ;
  assign n2347 = n2345 ^ x150 ;
  assign n2346 = n2345 ^ n2304 ;
  assign n2348 = n2347 ^ n2346 ;
  assign n2349 = n2309 & ~n2348 ;
  assign n2350 = n2349 ^ n2347 ;
  assign n2387 = n2386 ^ n1279 ;
  assign n2389 = n2387 ^ x149 ;
  assign n2388 = n2387 ^ n2345 ;
  assign n2390 = n2389 ^ n2388 ;
  assign n2391 = ~n2350 & n2390 ;
  assign n2392 = n2391 ^ n2389 ;
  assign n2398 = n2397 ^ n650 ;
  assign n2427 = n2426 ^ n2398 ;
  assign n2429 = n2427 ^ x148 ;
  assign n2428 = n2427 ^ n2387 ;
  assign n2430 = n2429 ^ n2428 ;
  assign n2431 = n2392 & ~n2430 ;
  assign n2432 = n2431 ^ n2429 ;
  assign n2435 = n2427 ^ x147 ;
  assign n2436 = n2432 & ~n2435 ;
  assign n2437 = n2436 ^ x147 ;
  assign n2475 = n2472 ^ n2437 ;
  assign n2476 = n2083 ^ n2076 ;
  assign n2477 = n2463 ^ n2444 ;
  assign n2478 = n1250 ^ x103 ;
  assign n2479 = n2478 ^ n2043 ;
  assign n2480 = n2479 ^ n2463 ;
  assign n2481 = n2480 ^ n2478 ;
  assign n2482 = n2477 & ~n2481 ;
  assign n2483 = n2482 ^ n2479 ;
  assign n2484 = n2483 ^ n2083 ;
  assign n2485 = n2476 & n2484 ;
  assign n2486 = n2485 ^ n2076 ;
  assign n2488 = n2486 ^ n649 ;
  assign n2487 = n2486 ^ n2466 ;
  assign n2489 = n2488 ^ n2487 ;
  assign n2490 = n2471 & n2489 ;
  assign n2491 = n2490 ^ n2488 ;
  assign n2492 = n2491 ^ n647 ;
  assign n2493 = n2492 ^ x146 ;
  assign n2494 = n2493 ^ n2437 ;
  assign n2495 = n2494 ^ n2492 ;
  assign n2496 = ~n2475 & n2495 ;
  assign n2497 = n2496 ^ n2493 ;
  assign n2501 = n2120 ^ n2083 ;
  assign n2500 = n2478 ^ n2120 ;
  assign n2502 = n2501 ^ n2500 ;
  assign n2503 = n2483 & n2502 ;
  assign n2504 = n2503 ^ n2501 ;
  assign n2505 = n2504 ^ n1505 ;
  assign n2506 = n2486 ^ n647 ;
  assign n2507 = ~n2491 & ~n2506 ;
  assign n2508 = n2507 ^ n647 ;
  assign n2509 = n2508 ^ n2113 ;
  assign n2510 = n2509 ^ n2120 ;
  assign n2511 = n2510 ^ n2508 ;
  assign n2512 = ~n2505 & n2511 ;
  assign n2513 = n2512 ^ n2509 ;
  assign n2514 = n2513 ^ n1414 ;
  assign n2516 = n2514 ^ x145 ;
  assign n2515 = n2514 ^ n2492 ;
  assign n2517 = n2516 ^ n2515 ;
  assign n2518 = ~n2497 & n2517 ;
  assign n2519 = n2518 ^ n2516 ;
  assign n2524 = n2120 ^ n1505 ;
  assign n2525 = ~n2504 & n2524 ;
  assign n2526 = n2525 ^ n2120 ;
  assign n2522 = n1506 ^ n1505 ;
  assign n2523 = n2522 ^ n2163 ;
  assign n2527 = n2526 ^ n2523 ;
  assign n2528 = ~n2193 & ~n2527 ;
  assign n2529 = n2528 ^ n1448 ;
  assign n2531 = n2529 ^ n1414 ;
  assign n2530 = n2529 ^ n2508 ;
  assign n2532 = n2531 ^ n2530 ;
  assign n2533 = ~n2513 & ~n2532 ;
  assign n2534 = n2533 ^ n2531 ;
  assign n2535 = n2534 ^ n646 ;
  assign n2537 = n2535 ^ x144 ;
  assign n2536 = n2535 ^ n2514 ;
  assign n2538 = n2537 ^ n2536 ;
  assign n2539 = n2519 & ~n2538 ;
  assign n2540 = n2539 ^ n2537 ;
  assign n2547 = n1509 ^ n1507 ;
  assign n2543 = n2526 ^ n2522 ;
  assign n2544 = n2526 ^ n2163 ;
  assign n2545 = n2543 & n2544 ;
  assign n2546 = n2545 ^ n2163 ;
  assign n2548 = n2547 ^ n2546 ;
  assign n2549 = n2548 ^ n2233 ;
  assign n2550 = n2198 & n2549 ;
  assign n2551 = n2550 ^ n2233 ;
  assign n2553 = n2551 ^ n646 ;
  assign n2552 = n2551 ^ n2529 ;
  assign n2554 = n2553 ^ n2552 ;
  assign n2555 = ~n2534 & n2554 ;
  assign n2556 = n2555 ^ n2553 ;
  assign n2557 = n2556 ^ n805 ;
  assign n2559 = n2557 ^ x159 ;
  assign n2558 = n2557 ^ n2535 ;
  assign n2560 = n2559 ^ n2558 ;
  assign n2561 = n2540 & ~n2560 ;
  assign n2562 = n2561 ^ n2559 ;
  assign n2579 = n1511 ^ n1510 ;
  assign n2571 = n2233 ^ n2198 ;
  assign n2572 = n2571 ^ n2546 ;
  assign n2573 = n2275 ^ n2240 ;
  assign n2574 = n2573 ^ n2547 ;
  assign n2575 = n2574 ^ n2573 ;
  assign n2576 = n2575 ^ n2546 ;
  assign n2577 = ~n2572 & ~n2576 ;
  assign n2578 = n2577 ^ n2574 ;
  assign n2580 = n2579 ^ n2578 ;
  assign n2581 = n2240 & n2580 ;
  assign n2582 = n2581 ^ n2275 ;
  assign n2584 = n2582 ^ n805 ;
  assign n2583 = n2582 ^ n2551 ;
  assign n2585 = n2584 ^ n2583 ;
  assign n2586 = n2556 & ~n2585 ;
  assign n2587 = n2586 ^ n2584 ;
  assign n2588 = n2587 ^ n893 ;
  assign n2590 = n2588 ^ x158 ;
  assign n2589 = n2588 ^ n2557 ;
  assign n2591 = n2590 ^ n2589 ;
  assign n2592 = ~n2562 & n2591 ;
  assign n2593 = n2592 ^ n2590 ;
  assign n2612 = n2283 ^ n2276 ;
  assign n2615 = n2579 ^ n2573 ;
  assign n2616 = n2578 & ~n2615 ;
  assign n2614 = n2573 ^ n2283 ;
  assign n2617 = n2616 ^ n2614 ;
  assign n2613 = n1513 ^ n1512 ;
  assign n2618 = n2617 ^ n2613 ;
  assign n2619 = n2612 & n2618 ;
  assign n2620 = n2619 ^ n2276 ;
  assign n2622 = n2620 ^ n893 ;
  assign n2621 = n2620 ^ n2582 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2624 = ~n2587 & n2623 ;
  assign n2625 = n2624 ^ n2622 ;
  assign n2626 = n2625 ^ n1588 ;
  assign n2628 = n2626 ^ x157 ;
  assign n2627 = n2626 ^ n2588 ;
  assign n2629 = n2628 ^ n2627 ;
  assign n2630 = n2593 & ~n2629 ;
  assign n2631 = n2630 ^ n2628 ;
  assign n2664 = n1515 ^ n1514 ;
  assign n2659 = n2325 ^ n2283 ;
  assign n2660 = n2659 ^ n2325 ;
  assign n2661 = n2660 ^ n2613 ;
  assign n2662 = n2617 & ~n2661 ;
  assign n2663 = n2662 ^ n2659 ;
  assign n2665 = n2664 ^ n2663 ;
  assign n2666 = n2324 & n2665 ;
  assign n2667 = n2666 ^ n1651 ;
  assign n2669 = n2667 ^ n1588 ;
  assign n2668 = n2667 ^ n2620 ;
  assign n2670 = n2669 ^ n2668 ;
  assign n2671 = ~n2625 & n2670 ;
  assign n2672 = n2671 ^ n2669 ;
  assign n2673 = n2672 ^ n1002 ;
  assign n2675 = n2673 ^ x156 ;
  assign n2674 = n2673 ^ n2626 ;
  assign n2676 = n2675 ^ n2674 ;
  assign n2677 = n2631 & ~n2676 ;
  assign n2678 = n2677 ^ n2675 ;
  assign n2703 = n2362 ^ n2355 ;
  assign n2709 = n1517 ^ n1516 ;
  assign n2705 = n2362 ^ n2325 ;
  assign n2704 = n2664 ^ n2362 ;
  assign n2706 = n2705 ^ n2704 ;
  assign n2707 = ~n2663 & ~n2706 ;
  assign n2708 = n2707 ^ n2705 ;
  assign n2710 = n2709 ^ n2708 ;
  assign n2711 = ~n2703 & ~n2710 ;
  assign n2712 = n2711 ^ n2355 ;
  assign n2714 = n2712 ^ n1002 ;
  assign n2713 = n2712 ^ n2667 ;
  assign n2715 = n2714 ^ n2713 ;
  assign n2716 = n2672 & n2715 ;
  assign n2717 = n2716 ^ n2714 ;
  assign n2718 = n2717 ^ n1023 ;
  assign n2720 = n2718 ^ x155 ;
  assign n2719 = n2718 ^ n2673 ;
  assign n2721 = n2720 ^ n2719 ;
  assign n2722 = n2678 & ~n2721 ;
  assign n2723 = n2722 ^ n2720 ;
  assign n2749 = n2411 ^ n2404 ;
  assign n2755 = n1519 ^ n1518 ;
  assign n2751 = n2411 ^ n2362 ;
  assign n2750 = n2709 ^ n2411 ;
  assign n2752 = n2751 ^ n2750 ;
  assign n2753 = n2708 & ~n2752 ;
  assign n2754 = n2753 ^ n2751 ;
  assign n2756 = n2755 ^ n2754 ;
  assign n2757 = ~n2749 & n2756 ;
  assign n2758 = n2757 ^ n2404 ;
  assign n2760 = n2758 ^ n1023 ;
  assign n2759 = n2758 ^ n2712 ;
  assign n2761 = n2760 ^ n2759 ;
  assign n2762 = n2717 & n2761 ;
  assign n2763 = n2762 ^ n2760 ;
  assign n2764 = n2763 ^ n1049 ;
  assign n2766 = n2764 ^ x154 ;
  assign n2765 = n2764 ^ n2718 ;
  assign n2767 = n2766 ^ n2765 ;
  assign n2768 = ~n2723 & n2767 ;
  assign n2769 = n2768 ^ n2766 ;
  assign n2770 = n2769 ^ x153 ;
  assign n2724 = n2723 ^ x154 ;
  assign n2679 = n2678 ^ x155 ;
  assign n2632 = n2631 ^ x156 ;
  assign n2594 = n2593 ^ x157 ;
  assign n1944 = n1905 & ~n1943 ;
  assign n1984 = n1983 ^ x142 ;
  assign n1985 = n1944 & n1984 ;
  assign n2025 = n2024 ^ x141 ;
  assign n2026 = n1985 & n2025 ;
  assign n2064 = n2063 ^ x140 ;
  assign n2065 = n2026 & n2064 ;
  assign n2105 = n2104 ^ x139 ;
  assign n2106 = ~n2065 & n2105 ;
  assign n2147 = n2146 ^ x138 ;
  assign n2148 = n2106 & ~n2147 ;
  assign n2185 = n2184 ^ x137 ;
  assign n2186 = n2148 & ~n2185 ;
  assign n2226 = n2225 ^ x136 ;
  assign n2227 = n2186 & ~n2226 ;
  assign n2268 = n2267 ^ x151 ;
  assign n2269 = n2227 & n2268 ;
  assign n2310 = n2309 ^ x150 ;
  assign n2311 = n2269 & ~n2310 ;
  assign n2351 = n2350 ^ x149 ;
  assign n2352 = ~n2311 & ~n2351 ;
  assign n2393 = n2392 ^ x148 ;
  assign n2394 = n2352 & n2393 ;
  assign n2433 = n2432 ^ x147 ;
  assign n2434 = n2394 & n2433 ;
  assign n2438 = n2437 ^ x146 ;
  assign n2473 = n2472 ^ n2438 ;
  assign n2474 = n2434 & ~n2473 ;
  assign n2498 = n2497 ^ x145 ;
  assign n2499 = n2474 & ~n2498 ;
  assign n2520 = n2519 ^ x144 ;
  assign n2521 = ~n2499 & ~n2520 ;
  assign n2541 = n2540 ^ x159 ;
  assign n2542 = ~n2521 & n2541 ;
  assign n2563 = n2562 ^ x158 ;
  assign n2595 = ~n2542 & n2563 ;
  assign n2633 = n2594 & ~n2595 ;
  assign n2680 = ~n2632 & ~n2633 ;
  assign n2725 = n2679 & ~n2680 ;
  assign n2748 = ~n2724 & n2725 ;
  assign n2771 = n2770 ^ n2748 ;
  assign n2788 = n2771 ^ n1795 ;
  assign n2726 = n2725 ^ n2724 ;
  assign n2743 = n2726 ^ n1733 ;
  assign n2681 = n2680 ^ n2679 ;
  assign n2698 = n2681 ^ n1676 ;
  assign n2634 = n2633 ^ n2632 ;
  assign n2654 = n2634 ^ n1620 ;
  assign n2564 = n2563 ^ n2542 ;
  assign n2597 = n1523 ^ n1183 ;
  assign n2598 = ~n2564 & n2597 ;
  assign n2599 = n2598 ^ n1571 ;
  assign n2596 = n2595 ^ n2594 ;
  assign n2608 = n2598 ^ n2596 ;
  assign n2609 = ~n2599 & ~n2608 ;
  assign n2610 = n2609 ^ n1571 ;
  assign n2655 = n2634 ^ n2610 ;
  assign n2656 = n2654 & n2655 ;
  assign n2657 = n2656 ^ n1620 ;
  assign n2699 = n2681 ^ n2657 ;
  assign n2700 = ~n2698 & ~n2699 ;
  assign n2701 = n2700 ^ n1676 ;
  assign n2744 = n2726 ^ n2701 ;
  assign n2745 = ~n2743 & n2744 ;
  assign n2746 = n2745 ^ n1733 ;
  assign n2789 = n2771 ^ n2746 ;
  assign n2790 = ~n2788 & ~n2789 ;
  assign n2791 = n2790 ^ n1795 ;
  assign n2792 = n2791 ^ n1853 ;
  assign n2809 = n1049 ^ x152 ;
  assign n2810 = n2809 ^ n2448 ;
  assign n2807 = n2758 ^ n1049 ;
  assign n2808 = ~n2763 & n2807 ;
  assign n2811 = n2810 ^ n2808 ;
  assign n2799 = n2454 ^ n1834 ;
  assign n2803 = n2755 ^ n2411 ;
  assign n2804 = ~n2754 & n2803 ;
  assign n2800 = n1521 ^ n1520 ;
  assign n2801 = n2800 ^ n2454 ;
  assign n2802 = n2801 ^ n2755 ;
  assign n2805 = n2804 ^ n2802 ;
  assign n2806 = ~n2799 & ~n2805 ;
  assign n2812 = n2811 ^ n2806 ;
  assign n2794 = n2764 ^ n2748 ;
  assign n2797 = n2769 & ~n2794 ;
  assign n2793 = n2769 ^ n2764 ;
  assign n2795 = n2794 ^ n2793 ;
  assign n2796 = x153 & ~n2795 ;
  assign n2798 = n2797 ^ n2796 ;
  assign n2813 = n2812 ^ n2798 ;
  assign n2830 = n2813 ^ n2791 ;
  assign n2831 = n2792 & n2830 ;
  assign n2832 = n2831 ^ n1853 ;
  assign n2851 = n2833 ^ n2832 ;
  assign n2852 = ~n2834 & n2851 ;
  assign n2854 = n2853 ^ n2852 ;
  assign n2873 = n1970 ^ n1929 ;
  assign n2855 = n1575 ^ n1528 ;
  assign n2872 = n2855 ^ n1970 ;
  assign n2874 = n2873 ^ n2872 ;
  assign n2875 = ~n2854 & ~n2874 ;
  assign n2876 = n2875 ^ n2873 ;
  assign n2895 = n2011 ^ n1970 ;
  assign n2877 = n1634 ^ n1576 ;
  assign n2894 = n2877 ^ n2011 ;
  assign n2896 = n2895 ^ n2894 ;
  assign n2897 = n2876 & ~n2896 ;
  assign n2898 = n2897 ^ n2895 ;
  assign n2917 = n2050 ^ n2011 ;
  assign n2899 = n1690 ^ n1635 ;
  assign n2916 = n2899 ^ n2050 ;
  assign n2918 = n2917 ^ n2916 ;
  assign n2919 = ~n2898 & n2918 ;
  assign n2920 = n2919 ^ n2917 ;
  assign n2943 = n2091 ^ n2050 ;
  assign n2921 = n1747 ^ n1691 ;
  assign n2942 = n2921 ^ n2091 ;
  assign n2944 = n2943 ^ n2942 ;
  assign n2945 = n2920 & n2944 ;
  assign n2946 = n2945 ^ n2943 ;
  assign n2947 = n1804 ^ n1748 ;
  assign n2962 = n2947 ^ n2091 ;
  assign n2963 = n2946 & n2962 ;
  assign n2961 = n2133 ^ n2091 ;
  assign n2964 = n2963 ^ n2961 ;
  assign n2960 = n1862 ^ n1805 ;
  assign n2982 = n2960 ^ n2133 ;
  assign n2983 = n2964 & n2982 ;
  assign n2985 = n2984 ^ n2983 ;
  assign n3002 = n2212 ^ n2176 ;
  assign n3003 = n3002 ^ n2212 ;
  assign n2981 = n1904 ^ n1863 ;
  assign n3004 = n3003 ^ n2981 ;
  assign n3005 = n2985 & ~n3004 ;
  assign n3006 = n3005 ^ n3002 ;
  assign n3008 = n3007 ^ n3006 ;
  assign n3009 = n2229 & n3008 ;
  assign n3010 = n3009 ^ n1782 ;
  assign n2986 = n2985 ^ n2981 ;
  assign n2987 = n2189 & ~n2986 ;
  assign n2988 = n2987 ^ n1721 ;
  assign n2997 = n2988 ^ n1126 ;
  assign n2965 = n2964 ^ n2960 ;
  assign n2966 = ~n2154 & n2965 ;
  assign n2967 = n2966 ^ n1663 ;
  assign n2976 = n2967 ^ n1644 ;
  assign n2948 = n2947 ^ n2946 ;
  assign n2949 = ~n2108 & n2948 ;
  assign n2950 = n2949 ^ n1606 ;
  assign n2955 = n2950 ^ n1586 ;
  assign n2922 = n2921 ^ n2920 ;
  assign n2923 = ~n2067 & n2922 ;
  assign n2924 = n2923 ^ n1556 ;
  assign n2937 = n2924 ^ n1537 ;
  assign n2900 = n2899 ^ n2898 ;
  assign n2901 = n2028 & ~n2900 ;
  assign n2902 = n2901 ^ n1493 ;
  assign n2911 = n2902 ^ n1060 ;
  assign n2878 = n2877 ^ n2876 ;
  assign n2879 = n1987 & n2878 ;
  assign n2880 = n2879 ^ n1460 ;
  assign n2889 = n2880 ^ n1033 ;
  assign n2856 = n2855 ^ n2854 ;
  assign n2857 = ~n1946 & ~n2856 ;
  assign n2858 = n2857 ^ n1427 ;
  assign n2867 = n2858 ^ n1408 ;
  assign n2835 = n2834 ^ n2832 ;
  assign n2836 = n1889 & ~n2835 ;
  assign n2837 = n2836 ^ n1394 ;
  assign n2814 = n2813 ^ n2792 ;
  assign n2815 = n1864 & ~n2814 ;
  assign n2816 = n2815 ^ n1360 ;
  assign n2825 = n2816 ^ n933 ;
  assign n2747 = n2746 ^ n1795 ;
  assign n2772 = n2771 ^ n2747 ;
  assign n2773 = n1812 & n2772 ;
  assign n2774 = n2773 ^ n1329 ;
  assign n2783 = n2774 ^ n929 ;
  assign n2702 = n2701 ^ n1733 ;
  assign n2727 = n2726 ^ n2702 ;
  assign n2728 = ~n1754 & n2727 ;
  assign n2729 = n2728 ^ n1298 ;
  assign n2738 = n2729 ^ n1274 ;
  assign n2658 = n2657 ^ n1676 ;
  assign n2682 = n2681 ^ n2658 ;
  assign n2683 = n1693 & ~n2682 ;
  assign n2684 = n2683 ^ n1245 ;
  assign n2693 = n2684 ^ n923 ;
  assign n2565 = n2564 ^ n1183 ;
  assign n2566 = ~n1523 & ~n2565 ;
  assign n2567 = n2566 ^ n1183 ;
  assign n2603 = ~n1182 & ~n2567 ;
  assign n2604 = n2603 ^ n917 ;
  assign n2600 = n2599 ^ n2596 ;
  assign n2601 = n1579 & ~n2600 ;
  assign n2602 = n2601 ^ n1251 ;
  assign n2638 = n2603 ^ n2602 ;
  assign n2639 = ~n2604 & n2638 ;
  assign n2640 = n2639 ^ n917 ;
  assign n2641 = n2640 ^ n920 ;
  assign n2611 = n2610 ^ n1620 ;
  assign n2635 = n2634 ^ n2611 ;
  assign n2636 = n1619 & ~n2635 ;
  assign n2637 = n2636 ^ n1256 ;
  assign n2650 = n2640 ^ n2637 ;
  assign n2651 = ~n2641 & n2650 ;
  assign n2652 = n2651 ^ n920 ;
  assign n2694 = n2684 ^ n2652 ;
  assign n2695 = n2693 & n2694 ;
  assign n2696 = n2695 ^ n923 ;
  assign n2739 = n2729 ^ n2696 ;
  assign n2740 = ~n2738 & n2739 ;
  assign n2741 = n2740 ^ n1274 ;
  assign n2784 = n2774 ^ n2741 ;
  assign n2785 = n2783 & n2784 ;
  assign n2786 = n2785 ^ n929 ;
  assign n2826 = n2816 ^ n2786 ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = n2827 ^ n933 ;
  assign n2846 = n2837 ^ n2828 ;
  assign n2847 = n2837 ^ n1374 ;
  assign n2848 = ~n2846 & n2847 ;
  assign n2849 = n2848 ^ n1374 ;
  assign n2868 = n2858 ^ n2849 ;
  assign n2869 = ~n2867 & n2868 ;
  assign n2870 = n2869 ^ n1408 ;
  assign n2890 = n2880 ^ n2870 ;
  assign n2891 = ~n2889 & ~n2890 ;
  assign n2892 = n2891 ^ n1033 ;
  assign n2912 = n2902 ^ n2892 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2914 = n2913 ^ n1060 ;
  assign n2938 = n2924 ^ n2914 ;
  assign n2939 = ~n2937 & ~n2938 ;
  assign n2940 = n2939 ^ n1537 ;
  assign n2956 = n2950 ^ n2940 ;
  assign n2957 = ~n2955 & n2956 ;
  assign n2958 = n2957 ^ n1586 ;
  assign n2977 = n2967 ^ n2958 ;
  assign n2978 = n2976 & n2977 ;
  assign n2979 = n2978 ^ n1644 ;
  assign n2998 = n2988 ^ n2979 ;
  assign n2999 = n2997 & n2998 ;
  assign n3000 = n2999 ^ n1126 ;
  assign n3019 = n3010 ^ n3000 ;
  assign n3022 = n3007 ^ n2212 ;
  assign n3023 = n3006 & n3022 ;
  assign n3024 = n3023 ^ n2212 ;
  assign n3020 = n1984 ^ n1944 ;
  assign n3021 = n3020 ^ n2254 ;
  assign n3025 = n3024 ^ n3021 ;
  assign n3026 = ~n2274 & ~n3025 ;
  assign n3027 = n3026 ^ n1841 ;
  assign n3028 = n3027 ^ n1763 ;
  assign n3029 = n3028 ^ n3000 ;
  assign n3030 = n3029 ^ n3027 ;
  assign n3031 = ~n3019 & n3030 ;
  assign n3032 = n3031 ^ n3028 ;
  assign n3045 = n3024 ^ n3020 ;
  assign n3046 = n2025 ^ n1985 ;
  assign n3047 = n3046 ^ n2254 ;
  assign n3048 = n3047 ^ n3024 ;
  assign n3049 = n3048 ^ n3046 ;
  assign n3050 = n3045 & n3049 ;
  assign n3051 = n3050 ^ n3047 ;
  assign n3052 = n3051 ^ n1872 ;
  assign n3053 = n2300 & ~n3052 ;
  assign n3054 = n3053 ^ n1872 ;
  assign n3056 = n3054 ^ n1191 ;
  assign n3055 = n3054 ^ n3027 ;
  assign n3057 = n3056 ^ n3055 ;
  assign n3058 = n3032 & n3057 ;
  assign n3059 = n3058 ^ n3056 ;
  assign n3060 = n3059 ^ n1211 ;
  assign n2941 = n2940 ^ n1586 ;
  assign n2951 = n2950 ^ n2941 ;
  assign n2605 = n2604 ^ n2602 ;
  assign n2568 = n2567 ^ n1182 ;
  assign n2569 = x167 & n2568 ;
  assign n2607 = n2605 ^ n2569 ;
  assign n2642 = n2641 ^ n2637 ;
  assign n2643 = n2642 ^ x166 ;
  assign n2644 = n2643 ^ n2605 ;
  assign n2645 = n2644 ^ n2642 ;
  assign n2646 = ~n2607 & n2645 ;
  assign n2647 = n2646 ^ n2643 ;
  assign n2653 = n2652 ^ n923 ;
  assign n2685 = n2684 ^ n2653 ;
  assign n2687 = n2685 ^ x165 ;
  assign n2686 = n2685 ^ n2642 ;
  assign n2688 = n2687 ^ n2686 ;
  assign n2689 = n2647 & ~n2688 ;
  assign n2690 = n2689 ^ n2687 ;
  assign n2697 = n2696 ^ n1274 ;
  assign n2730 = n2729 ^ n2697 ;
  assign n2732 = n2730 ^ x164 ;
  assign n2731 = n2730 ^ n2685 ;
  assign n2733 = n2732 ^ n2731 ;
  assign n2734 = ~n2690 & n2733 ;
  assign n2735 = n2734 ^ n2732 ;
  assign n2742 = n2741 ^ n929 ;
  assign n2775 = n2774 ^ n2742 ;
  assign n2777 = n2775 ^ x163 ;
  assign n2776 = n2775 ^ n2730 ;
  assign n2778 = n2777 ^ n2776 ;
  assign n2779 = ~n2735 & n2778 ;
  assign n2780 = n2779 ^ n2777 ;
  assign n2787 = n2786 ^ n933 ;
  assign n2817 = n2816 ^ n2787 ;
  assign n2819 = n2817 ^ x162 ;
  assign n2818 = n2817 ^ n2775 ;
  assign n2820 = n2819 ^ n2818 ;
  assign n2821 = n2780 & ~n2820 ;
  assign n2822 = n2821 ^ n2819 ;
  assign n2829 = n2828 ^ n1374 ;
  assign n2838 = n2837 ^ n2829 ;
  assign n2840 = n2838 ^ x161 ;
  assign n2839 = n2838 ^ n2817 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2842 = n2822 & ~n2841 ;
  assign n2843 = n2842 ^ n2840 ;
  assign n2850 = n2849 ^ n1408 ;
  assign n2859 = n2858 ^ n2850 ;
  assign n2861 = n2859 ^ x160 ;
  assign n2860 = n2859 ^ n2838 ;
  assign n2862 = n2861 ^ n2860 ;
  assign n2863 = n2843 & ~n2862 ;
  assign n2864 = n2863 ^ n2861 ;
  assign n2871 = n2870 ^ n1033 ;
  assign n2881 = n2880 ^ n2871 ;
  assign n2883 = n2881 ^ x175 ;
  assign n2882 = n2881 ^ n2859 ;
  assign n2884 = n2883 ^ n2882 ;
  assign n2885 = ~n2864 & n2884 ;
  assign n2886 = n2885 ^ n2883 ;
  assign n2893 = n2892 ^ n1060 ;
  assign n2903 = n2902 ^ n2893 ;
  assign n2905 = n2903 ^ x174 ;
  assign n2904 = n2903 ^ n2881 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n2907 = ~n2886 & n2906 ;
  assign n2908 = n2907 ^ n2905 ;
  assign n2915 = n2914 ^ n1537 ;
  assign n2925 = n2924 ^ n2915 ;
  assign n2927 = n2925 ^ x173 ;
  assign n2926 = n2925 ^ n2903 ;
  assign n2928 = n2927 ^ n2926 ;
  assign n2929 = n2908 & ~n2928 ;
  assign n2930 = n2929 ^ n2927 ;
  assign n2933 = n2925 ^ x172 ;
  assign n2934 = ~n2930 & n2933 ;
  assign n2935 = n2934 ^ x172 ;
  assign n2954 = n2951 ^ n2935 ;
  assign n2959 = n2958 ^ n1644 ;
  assign n2968 = n2967 ^ n2959 ;
  assign n2969 = n2968 ^ x171 ;
  assign n2970 = n2969 ^ n2935 ;
  assign n2971 = n2970 ^ n2968 ;
  assign n2972 = n2954 & n2971 ;
  assign n2973 = n2972 ^ n2969 ;
  assign n2980 = n2979 ^ n1126 ;
  assign n2989 = n2988 ^ n2980 ;
  assign n2991 = n2989 ^ x170 ;
  assign n2990 = n2989 ^ n2968 ;
  assign n2992 = n2991 ^ n2990 ;
  assign n2993 = ~n2973 & n2992 ;
  assign n2994 = n2993 ^ n2991 ;
  assign n3001 = n3000 ^ n1763 ;
  assign n3011 = n3010 ^ n3001 ;
  assign n3013 = n3011 ^ x169 ;
  assign n3012 = n3011 ^ n2989 ;
  assign n3014 = n3013 ^ n3012 ;
  assign n3015 = n2994 & ~n3014 ;
  assign n3016 = n3015 ^ n3013 ;
  assign n3033 = n3032 ^ n1191 ;
  assign n3035 = n3033 ^ x168 ;
  assign n3034 = n3033 ^ n3011 ;
  assign n3036 = n3035 ^ n3034 ;
  assign n3037 = ~n3016 & n3036 ;
  assign n3038 = n3037 ^ n3035 ;
  assign n3041 = n3033 ^ x183 ;
  assign n3042 = ~n3038 & n3041 ;
  assign n3043 = n3042 ^ x183 ;
  assign n3063 = n3060 ^ n3043 ;
  assign n3069 = n2064 ^ n2026 ;
  assign n3067 = n3046 ^ n2337 ;
  assign n3064 = n2300 ^ n1872 ;
  assign n3065 = n3064 ^ n3046 ;
  assign n3066 = ~n3051 & n3065 ;
  assign n3068 = n3067 ^ n3066 ;
  assign n3070 = n3069 ^ n3068 ;
  assign n3071 = n2375 & ~n3070 ;
  assign n3072 = n3071 ^ n1916 ;
  assign n3074 = n3072 ^ n1211 ;
  assign n3073 = n3072 ^ n3054 ;
  assign n3075 = n3074 ^ n3073 ;
  assign n3076 = ~n3059 & n3075 ;
  assign n3077 = n3076 ^ n3074 ;
  assign n3078 = n3077 ^ n1913 ;
  assign n3079 = n3078 ^ x182 ;
  assign n3080 = n3079 ^ n3043 ;
  assign n3081 = n3080 ^ n3078 ;
  assign n3082 = n3063 & n3081 ;
  assign n3083 = n3082 ^ n3079 ;
  assign n3094 = n3072 ^ n1913 ;
  assign n3095 = ~n3077 & ~n3094 ;
  assign n3096 = n3095 ^ n1913 ;
  assign n3097 = n3096 ^ n1286 ;
  assign n3088 = n3069 ^ n2337 ;
  assign n3089 = n3068 & n3088 ;
  assign n3087 = n2379 ^ n2337 ;
  assign n3090 = n3089 ^ n3087 ;
  assign n3086 = n2105 ^ n2065 ;
  assign n3091 = n3090 ^ n3086 ;
  assign n3092 = ~n2400 & ~n3091 ;
  assign n3093 = n3092 ^ n1956 ;
  assign n3098 = n3097 ^ n3093 ;
  assign n3100 = n3098 ^ x181 ;
  assign n3099 = n3098 ^ n3078 ;
  assign n3101 = n3100 ^ n3099 ;
  assign n3102 = ~n3083 & n3101 ;
  assign n3103 = n3102 ^ n3100 ;
  assign n3114 = n3096 ^ n3093 ;
  assign n3115 = ~n3097 & ~n3114 ;
  assign n3116 = n3115 ^ n1286 ;
  assign n3117 = n3116 ^ n1315 ;
  assign n3109 = n2424 ^ n2379 ;
  assign n3107 = n3086 ^ n2379 ;
  assign n3108 = n3090 & n3107 ;
  assign n3110 = n3109 ^ n3108 ;
  assign n3106 = n2147 ^ n2106 ;
  assign n3111 = n3110 ^ n3106 ;
  assign n3112 = n2442 & n3111 ;
  assign n3113 = n3112 ^ n1997 ;
  assign n3118 = n3117 ^ n3113 ;
  assign n3120 = n3118 ^ x180 ;
  assign n3119 = n3118 ^ n3098 ;
  assign n3121 = n3120 ^ n3119 ;
  assign n3122 = n3103 & ~n3121 ;
  assign n3123 = n3122 ^ n3120 ;
  assign n3124 = n3123 ^ x179 ;
  assign n2570 = n2569 ^ x166 ;
  assign n2606 = n2605 ^ n2570 ;
  assign n2648 = n2647 ^ x165 ;
  assign n2649 = n2606 & ~n2648 ;
  assign n2691 = n2690 ^ x164 ;
  assign n2692 = ~n2649 & ~n2691 ;
  assign n2736 = n2735 ^ x163 ;
  assign n2737 = ~n2692 & n2736 ;
  assign n2781 = n2780 ^ x162 ;
  assign n2782 = ~n2737 & n2781 ;
  assign n2823 = n2822 ^ x161 ;
  assign n2824 = ~n2782 & ~n2823 ;
  assign n2844 = n2843 ^ x160 ;
  assign n2845 = n2824 & ~n2844 ;
  assign n2865 = n2864 ^ x175 ;
  assign n2866 = n2845 & n2865 ;
  assign n2887 = n2886 ^ x174 ;
  assign n2888 = ~n2866 & ~n2887 ;
  assign n2909 = n2908 ^ x173 ;
  assign n2910 = n2888 & n2909 ;
  assign n2931 = n2930 ^ x172 ;
  assign n2932 = ~n2910 & n2931 ;
  assign n2936 = n2935 ^ x171 ;
  assign n2952 = n2951 ^ n2936 ;
  assign n2953 = n2932 & ~n2952 ;
  assign n2974 = n2973 ^ x170 ;
  assign n2975 = n2953 & n2974 ;
  assign n2995 = n2994 ^ x169 ;
  assign n2996 = ~n2975 & n2995 ;
  assign n3017 = n3016 ^ x168 ;
  assign n3018 = n2996 & ~n3017 ;
  assign n3039 = n3038 ^ x183 ;
  assign n3040 = n3018 & ~n3039 ;
  assign n3044 = n3043 ^ x182 ;
  assign n3061 = n3060 ^ n3044 ;
  assign n3062 = n3040 & n3061 ;
  assign n3084 = n3083 ^ x181 ;
  assign n3085 = n3062 & ~n3084 ;
  assign n3104 = n3103 ^ x180 ;
  assign n3105 = ~n3085 & ~n3104 ;
  assign n3125 = n3124 ^ n3105 ;
  assign n3126 = n3125 ^ n2597 ;
  assign n3127 = ~n2564 & ~n3126 ;
  assign n3128 = n3127 ^ n2597 ;
  assign n3161 = n3128 ^ n1183 ;
  assign n3162 = x199 & ~n3161 ;
  assign n3138 = n3116 ^ n3113 ;
  assign n3144 = n2185 ^ n2148 ;
  assign n3139 = n2464 ^ n2424 ;
  assign n3140 = n3139 ^ n2464 ;
  assign n3141 = n3140 ^ n3106 ;
  assign n3142 = ~n3110 & ~n3141 ;
  assign n3143 = n3142 ^ n3139 ;
  assign n3145 = n3144 ^ n3143 ;
  assign n3146 = ~n2477 & n3145 ;
  assign n3147 = n3146 ^ n2043 ;
  assign n3148 = n3147 ^ n1315 ;
  assign n3149 = n3148 ^ n3113 ;
  assign n3150 = n3149 ^ n3147 ;
  assign n3151 = n3138 & ~n3150 ;
  assign n3152 = n3151 ^ n3148 ;
  assign n3153 = n3152 ^ n1348 ;
  assign n3135 = n3118 ^ x179 ;
  assign n3136 = ~n3123 & n3135 ;
  assign n3137 = n3136 ^ x179 ;
  assign n3154 = n3153 ^ n3137 ;
  assign n3155 = n3154 ^ x178 ;
  assign n3134 = n3105 & n3124 ;
  assign n3156 = n3155 ^ n3134 ;
  assign n3131 = n2597 ^ n2564 ;
  assign n3132 = n3125 & ~n3131 ;
  assign n3133 = n3132 ^ n2600 ;
  assign n3157 = n3156 ^ n3133 ;
  assign n3158 = n2608 & ~n3157 ;
  assign n3159 = n3158 ^ n1571 ;
  assign n3129 = ~n1183 & n3128 ;
  assign n3130 = n3129 ^ n1251 ;
  assign n3160 = n3159 ^ n3130 ;
  assign n3163 = n3162 ^ n3160 ;
  assign n3184 = n3147 ^ n1348 ;
  assign n3185 = n3152 & ~n3184 ;
  assign n3186 = n3185 ^ n1348 ;
  assign n3187 = n3186 ^ n2076 ;
  assign n3180 = n2226 ^ n2186 ;
  assign n3176 = n2484 ^ n2464 ;
  assign n3175 = n3144 ^ n2484 ;
  assign n3177 = n3176 ^ n3175 ;
  assign n3178 = ~n3143 & n3177 ;
  assign n3179 = n3178 ^ n3176 ;
  assign n3181 = n3180 ^ n3179 ;
  assign n3182 = ~n2483 & n3181 ;
  assign n3183 = n3182 ^ n2083 ;
  assign n3188 = n3187 ^ n3183 ;
  assign n3189 = n3188 ^ x178 ;
  assign n3190 = n3189 ^ n3137 ;
  assign n3191 = n3190 ^ n3188 ;
  assign n3192 = ~n3154 & n3191 ;
  assign n3193 = n3192 ^ n3189 ;
  assign n3194 = n3193 ^ x177 ;
  assign n3174 = n3134 & n3155 ;
  assign n3195 = n3194 ^ n3174 ;
  assign n3169 = n3156 ^ n3132 ;
  assign n3170 = n3156 ^ n2600 ;
  assign n3171 = ~n3169 & ~n3170 ;
  assign n3172 = n3171 ^ n2600 ;
  assign n3173 = n3172 ^ n2635 ;
  assign n3196 = n3195 ^ n3173 ;
  assign n3197 = ~n2655 & ~n3196 ;
  assign n3198 = n3197 ^ n1620 ;
  assign n3164 = n3159 ^ n3129 ;
  assign n3165 = n3159 ^ n1251 ;
  assign n3166 = n3164 & n3165 ;
  assign n3167 = n3166 ^ n1251 ;
  assign n3168 = n3167 ^ n1256 ;
  assign n3199 = n3198 ^ n3168 ;
  assign n3200 = n3199 ^ x198 ;
  assign n3201 = n3200 ^ n3160 ;
  assign n3202 = n3201 ^ n3199 ;
  assign n3203 = ~n3163 & n3202 ;
  assign n3204 = n3203 ^ n3200 ;
  assign n3232 = n3195 ^ n3172 ;
  assign n3233 = n3195 ^ n2635 ;
  assign n3234 = ~n3232 & n3233 ;
  assign n3235 = n3234 ^ n2635 ;
  assign n3236 = n3235 ^ n2682 ;
  assign n3220 = n3186 ^ n3183 ;
  assign n3221 = n3187 & ~n3220 ;
  assign n3222 = n3221 ^ n2076 ;
  assign n3223 = n3222 ^ n2113 ;
  assign n3211 = n2505 ^ n2120 ;
  assign n3213 = n3180 ^ n2484 ;
  assign n3214 = ~n3179 & ~n3213 ;
  assign n3215 = n3214 ^ n2484 ;
  assign n3212 = n2268 ^ n2227 ;
  assign n3216 = n3215 ^ n3212 ;
  assign n3217 = n3216 ^ n2505 ;
  assign n3218 = ~n3211 & ~n3217 ;
  assign n3219 = n3218 ^ n2120 ;
  assign n3224 = n3223 ^ n3219 ;
  assign n3226 = n3224 ^ x177 ;
  assign n3225 = n3224 ^ n3188 ;
  assign n3227 = n3226 ^ n3225 ;
  assign n3228 = n3193 & ~n3227 ;
  assign n3229 = n3228 ^ n3226 ;
  assign n3230 = n3229 ^ x176 ;
  assign n3210 = n3174 & ~n3194 ;
  assign n3231 = n3230 ^ n3210 ;
  assign n3237 = n3236 ^ n3231 ;
  assign n3238 = n2699 & n3237 ;
  assign n3239 = n3238 ^ n1676 ;
  assign n3205 = n3198 ^ n3167 ;
  assign n3206 = n3198 ^ n1256 ;
  assign n3207 = n3205 & n3206 ;
  assign n3208 = n3207 ^ n1256 ;
  assign n3209 = n3208 ^ n1245 ;
  assign n3240 = n3239 ^ n3209 ;
  assign n3242 = n3240 ^ x197 ;
  assign n3241 = n3240 ^ n3199 ;
  assign n3243 = n3242 ^ n3241 ;
  assign n3244 = n3204 & ~n3243 ;
  assign n3245 = n3244 ^ n3242 ;
  assign n3257 = n3222 ^ n3219 ;
  assign n3258 = n2310 ^ n2269 ;
  assign n3259 = n3258 ^ n2505 ;
  assign n3260 = n3259 ^ n3215 ;
  assign n3261 = n3260 ^ n3258 ;
  assign n3262 = ~n3216 & ~n3261 ;
  assign n3263 = n3262 ^ n3259 ;
  assign n3264 = n3263 ^ n2163 ;
  assign n3265 = ~n2543 & ~n3264 ;
  assign n3266 = n3265 ^ n2163 ;
  assign n3267 = n3266 ^ n2113 ;
  assign n3268 = n3267 ^ n3219 ;
  assign n3269 = n3268 ^ n3266 ;
  assign n3270 = n3257 & n3269 ;
  assign n3271 = n3270 ^ n3267 ;
  assign n3272 = n3271 ^ n1448 ;
  assign n3274 = n3272 ^ x176 ;
  assign n3273 = n3272 ^ n3224 ;
  assign n3275 = n3274 ^ n3273 ;
  assign n3276 = n3229 & ~n3275 ;
  assign n3277 = n3276 ^ n3274 ;
  assign n3278 = n3277 ^ x191 ;
  assign n3256 = ~n3210 & n3230 ;
  assign n3279 = n3278 ^ n3256 ;
  assign n3251 = n3235 ^ n3231 ;
  assign n3252 = n3231 ^ n2682 ;
  assign n3253 = n3251 & ~n3252 ;
  assign n3254 = n3253 ^ n2682 ;
  assign n3255 = n3254 ^ n2727 ;
  assign n3280 = n3279 ^ n3255 ;
  assign n3281 = ~n2744 & n3280 ;
  assign n3282 = n3281 ^ n1733 ;
  assign n3246 = n3239 ^ n3208 ;
  assign n3247 = n3239 ^ n1245 ;
  assign n3248 = n3246 & n3247 ;
  assign n3249 = n3248 ^ n1245 ;
  assign n3250 = n3249 ^ n1298 ;
  assign n3283 = n3282 ^ n3250 ;
  assign n3285 = n3283 ^ x196 ;
  assign n3284 = n3283 ^ n3240 ;
  assign n3286 = n3285 ^ n3284 ;
  assign n3287 = ~n3245 & n3286 ;
  assign n3288 = n3287 ^ n3285 ;
  assign n3318 = n3279 ^ n3254 ;
  assign n3319 = n3279 ^ n2727 ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = n3320 ^ n2727 ;
  assign n3322 = n3321 ^ n2772 ;
  assign n3301 = n2351 ^ n2311 ;
  assign n3295 = n2571 ^ n2548 ;
  assign n3297 = n3295 ^ n2527 ;
  assign n3296 = n3295 ^ n3258 ;
  assign n3298 = n3297 ^ n3296 ;
  assign n3299 = ~n3263 & n3298 ;
  assign n3300 = n3299 ^ n3297 ;
  assign n3302 = n3301 ^ n3300 ;
  assign n3303 = ~n2548 & ~n3302 ;
  assign n3304 = n3303 ^ n2571 ;
  assign n3306 = n3304 ^ n1448 ;
  assign n3305 = n3304 ^ n3266 ;
  assign n3307 = n3306 ^ n3305 ;
  assign n3308 = ~n3271 & ~n3307 ;
  assign n3309 = n3308 ^ n3306 ;
  assign n3310 = n3309 ^ n2233 ;
  assign n3312 = n3310 ^ x191 ;
  assign n3311 = n3310 ^ n3272 ;
  assign n3313 = n3312 ^ n3311 ;
  assign n3314 = n3277 & ~n3313 ;
  assign n3315 = n3314 ^ n3312 ;
  assign n3316 = n3315 ^ x190 ;
  assign n3294 = n3256 & n3278 ;
  assign n3317 = n3316 ^ n3294 ;
  assign n3323 = n3322 ^ n3317 ;
  assign n3324 = n2789 & ~n3323 ;
  assign n3325 = n3324 ^ n1795 ;
  assign n3289 = n3282 ^ n3249 ;
  assign n3290 = n3282 ^ n1298 ;
  assign n3291 = ~n3289 & ~n3290 ;
  assign n3292 = n3291 ^ n1298 ;
  assign n3293 = n3292 ^ n1329 ;
  assign n3326 = n3325 ^ n3293 ;
  assign n3328 = n3326 ^ x195 ;
  assign n3327 = n3326 ^ n3283 ;
  assign n3329 = n3328 ^ n3327 ;
  assign n3330 = ~n3288 & n3329 ;
  assign n3331 = n3330 ^ n3328 ;
  assign n3346 = n2580 ^ n2573 ;
  assign n3349 = n3301 ^ n3295 ;
  assign n3350 = n3300 & n3349 ;
  assign n3348 = n3295 ^ n2580 ;
  assign n3351 = n3350 ^ n3348 ;
  assign n3347 = n2393 ^ n2352 ;
  assign n3352 = n3351 ^ n3347 ;
  assign n3353 = ~n3346 & n3352 ;
  assign n3354 = n3353 ^ n2573 ;
  assign n3342 = n3304 ^ n2233 ;
  assign n3343 = n3309 & n3342 ;
  assign n3344 = n3343 ^ n2233 ;
  assign n3345 = n3344 ^ n2275 ;
  assign n3355 = n3354 ^ n3345 ;
  assign n3357 = n3355 ^ x190 ;
  assign n3356 = n3355 ^ n3310 ;
  assign n3358 = n3357 ^ n3356 ;
  assign n3359 = n3315 & ~n3358 ;
  assign n3360 = n3359 ^ n3357 ;
  assign n3361 = n3360 ^ x189 ;
  assign n3341 = n3294 & n3316 ;
  assign n3362 = n3361 ^ n3341 ;
  assign n3337 = n3321 ^ n3317 ;
  assign n3338 = n3322 & n3337 ;
  assign n3339 = n3338 ^ n2772 ;
  assign n3340 = n3339 ^ n2814 ;
  assign n3363 = n3362 ^ n3340 ;
  assign n3364 = ~n2830 & ~n3363 ;
  assign n3365 = n3364 ^ n1853 ;
  assign n3332 = n3325 ^ n3292 ;
  assign n3333 = n3325 ^ n1329 ;
  assign n3334 = ~n3332 & n3333 ;
  assign n3335 = n3334 ^ n1329 ;
  assign n3336 = n3335 ^ n1360 ;
  assign n3366 = n3365 ^ n3336 ;
  assign n3368 = n3366 ^ x194 ;
  assign n3367 = n3366 ^ n3326 ;
  assign n3369 = n3368 ^ n3367 ;
  assign n3370 = ~n3331 & n3369 ;
  assign n3371 = n3370 ^ n3368 ;
  assign n3377 = n2832 ^ n1528 ;
  assign n3401 = n3362 ^ n3339 ;
  assign n3402 = n3362 ^ n2814 ;
  assign n3403 = ~n3401 & ~n3402 ;
  assign n3404 = n3403 ^ n2814 ;
  assign n3405 = n3404 ^ n2835 ;
  assign n3395 = n3355 ^ x189 ;
  assign n3396 = ~n3360 & n3395 ;
  assign n3397 = n3396 ^ x189 ;
  assign n3398 = n3397 ^ x188 ;
  assign n3384 = n2618 ^ n2283 ;
  assign n3390 = n2433 ^ n2394 ;
  assign n3385 = n2618 ^ n2580 ;
  assign n3386 = n3385 ^ n2618 ;
  assign n3387 = n3386 ^ n3347 ;
  assign n3388 = ~n3351 & ~n3387 ;
  assign n3389 = n3388 ^ n3385 ;
  assign n3391 = n3390 ^ n3389 ;
  assign n3392 = ~n3384 & ~n3391 ;
  assign n3393 = n3392 ^ n2283 ;
  assign n3379 = n3354 ^ n3344 ;
  assign n3380 = n3354 ^ n2275 ;
  assign n3381 = n3379 & n3380 ;
  assign n3382 = n3381 ^ n2275 ;
  assign n3383 = n3382 ^ n2276 ;
  assign n3394 = n3393 ^ n3383 ;
  assign n3399 = n3398 ^ n3394 ;
  assign n3378 = n3341 & ~n3361 ;
  assign n3400 = n3399 ^ n3378 ;
  assign n3406 = n3405 ^ n3400 ;
  assign n3407 = n3377 & n3406 ;
  assign n3408 = n3407 ^ n2833 ;
  assign n3372 = n3365 ^ n3335 ;
  assign n3373 = n3365 ^ n1360 ;
  assign n3374 = ~n3372 & n3373 ;
  assign n3375 = n3374 ^ n1360 ;
  assign n3376 = n3375 ^ n1394 ;
  assign n3409 = n3408 ^ n3376 ;
  assign n3411 = n3409 ^ x193 ;
  assign n3410 = n3409 ^ n3366 ;
  assign n3412 = n3411 ^ n3410 ;
  assign n3413 = ~n3371 & n3412 ;
  assign n3414 = n3413 ^ n3411 ;
  assign n3415 = n3414 ^ x192 ;
  assign n3416 = n3161 ^ x199 ;
  assign n3417 = n3162 ^ x198 ;
  assign n3418 = n3417 ^ n3160 ;
  assign n3419 = n3416 & ~n3418 ;
  assign n3420 = n3204 ^ x197 ;
  assign n3421 = ~n3419 & ~n3420 ;
  assign n3422 = n3245 ^ x196 ;
  assign n3423 = n3421 & n3422 ;
  assign n3424 = n3288 ^ x195 ;
  assign n3425 = ~n3423 & ~n3424 ;
  assign n3426 = n3331 ^ x194 ;
  assign n3427 = ~n3425 & n3426 ;
  assign n3428 = n3371 ^ x193 ;
  assign n3429 = n3427 & n3428 ;
  assign n3996 = n3415 & n3429 ;
  assign n3631 = n3408 ^ n3375 ;
  assign n3632 = n3408 ^ n1394 ;
  assign n3633 = n3631 & n3632 ;
  assign n3634 = n3633 ^ n1394 ;
  assign n3824 = n3634 ^ n1427 ;
  assign n3635 = n2856 ^ n1929 ;
  assign n3437 = n3404 ^ n3400 ;
  assign n3438 = n3400 ^ n2835 ;
  assign n3439 = n3437 & ~n3438 ;
  assign n3440 = n3439 ^ n2835 ;
  assign n3636 = n3440 ^ n2856 ;
  assign n3442 = n3397 ^ n3394 ;
  assign n3448 = n2665 ^ n2325 ;
  assign n3454 = n2473 ^ n2434 ;
  assign n3450 = n2665 ^ n2618 ;
  assign n3449 = n3390 ^ n2665 ;
  assign n3451 = n3450 ^ n3449 ;
  assign n3452 = n3389 & ~n3451 ;
  assign n3453 = n3452 ^ n3450 ;
  assign n3455 = n3454 ^ n3453 ;
  assign n3456 = n3448 & n3455 ;
  assign n3457 = n3456 ^ n2325 ;
  assign n3443 = n3393 ^ n3382 ;
  assign n3444 = n3393 ^ n2276 ;
  assign n3445 = ~n3443 & n3444 ;
  assign n3446 = n3445 ^ n2276 ;
  assign n3447 = n3446 ^ n1651 ;
  assign n3458 = n3457 ^ n3447 ;
  assign n3459 = n3458 ^ x188 ;
  assign n3460 = n3459 ^ n3394 ;
  assign n3461 = n3460 ^ n3458 ;
  assign n3462 = n3442 & ~n3461 ;
  assign n3463 = n3462 ^ n3459 ;
  assign n3464 = n3463 ^ x187 ;
  assign n3441 = ~n3378 & ~n3399 ;
  assign n3465 = n3464 ^ n3441 ;
  assign n3637 = n3636 ^ n3465 ;
  assign n3638 = n3635 & ~n3637 ;
  assign n3639 = n3638 ^ n1929 ;
  assign n3825 = n3824 ^ n3639 ;
  assign n3827 = n3825 ^ x192 ;
  assign n3826 = n3825 ^ n3409 ;
  assign n3828 = n3827 ^ n3826 ;
  assign n3829 = ~n3414 & n3828 ;
  assign n3830 = n3829 ^ n3827 ;
  assign n3997 = n3830 ^ x207 ;
  assign n3998 = n3996 & n3997 ;
  assign n3640 = n3639 ^ n3634 ;
  assign n3641 = n3639 ^ n1427 ;
  assign n3642 = ~n3640 & ~n3641 ;
  assign n3643 = n3642 ^ n1427 ;
  assign n3831 = n3643 ^ n1460 ;
  assign n3644 = n2878 ^ n1970 ;
  assign n3493 = n3441 & ~n3464 ;
  assign n3476 = n2710 ^ n2362 ;
  assign n3482 = n2498 ^ n2474 ;
  assign n3478 = n2710 ^ n2665 ;
  assign n3477 = n3454 ^ n2710 ;
  assign n3479 = n3478 ^ n3477 ;
  assign n3480 = n3453 & n3479 ;
  assign n3481 = n3480 ^ n3478 ;
  assign n3483 = n3482 ^ n3481 ;
  assign n3484 = ~n3476 & ~n3483 ;
  assign n3485 = n3484 ^ n2362 ;
  assign n3471 = n3457 ^ n3446 ;
  assign n3472 = n3457 ^ n1651 ;
  assign n3473 = n3471 & n3472 ;
  assign n3474 = n3473 ^ n1651 ;
  assign n3475 = n3474 ^ n2355 ;
  assign n3486 = n3485 ^ n3475 ;
  assign n3488 = n3486 ^ x187 ;
  assign n3487 = n3486 ^ n3458 ;
  assign n3489 = n3488 ^ n3487 ;
  assign n3490 = n3463 & ~n3489 ;
  assign n3491 = n3490 ^ n3488 ;
  assign n3492 = n3491 ^ x186 ;
  assign n3494 = n3493 ^ n3492 ;
  assign n3466 = n3465 ^ n3440 ;
  assign n3467 = n3465 ^ n2856 ;
  assign n3468 = ~n3466 & n3467 ;
  assign n3469 = n3468 ^ n2856 ;
  assign n3470 = n3469 ^ n2878 ;
  assign n3645 = n3494 ^ n3470 ;
  assign n3646 = ~n3644 & n3645 ;
  assign n3647 = n3646 ^ n1970 ;
  assign n3832 = n3831 ^ n3647 ;
  assign n3834 = n3832 ^ x207 ;
  assign n3833 = n3832 ^ n3825 ;
  assign n3835 = n3834 ^ n3833 ;
  assign n3836 = ~n3830 & n3835 ;
  assign n3837 = n3836 ^ n3834 ;
  assign n3999 = n3837 ^ x206 ;
  assign n4000 = ~n3998 & ~n3999 ;
  assign n3648 = n3647 ^ n3643 ;
  assign n3649 = n3647 ^ n1460 ;
  assign n3650 = n3648 & n3649 ;
  assign n3651 = n3650 ^ n1460 ;
  assign n3838 = n3651 ^ n1493 ;
  assign n3652 = n2900 ^ n2011 ;
  assign n3495 = n3494 ^ n3469 ;
  assign n3496 = ~n3470 & ~n3495 ;
  assign n3497 = n3496 ^ n2878 ;
  assign n3653 = n3497 ^ n2900 ;
  assign n3520 = ~n3492 & n3493 ;
  assign n3503 = n2756 ^ n2411 ;
  assign n3509 = n2520 ^ n2499 ;
  assign n3505 = n2756 ^ n2710 ;
  assign n3504 = n3482 ^ n2756 ;
  assign n3506 = n3505 ^ n3504 ;
  assign n3507 = ~n3481 & ~n3506 ;
  assign n3508 = n3507 ^ n3505 ;
  assign n3510 = n3509 ^ n3508 ;
  assign n3511 = n3503 & ~n3510 ;
  assign n3512 = n3511 ^ n2411 ;
  assign n3498 = n3485 ^ n3474 ;
  assign n3499 = n3485 ^ n2355 ;
  assign n3500 = ~n3498 & ~n3499 ;
  assign n3501 = n3500 ^ n2355 ;
  assign n3502 = n3501 ^ n2404 ;
  assign n3513 = n3512 ^ n3502 ;
  assign n3515 = n3513 ^ x186 ;
  assign n3514 = n3513 ^ n3486 ;
  assign n3516 = n3515 ^ n3514 ;
  assign n3517 = n3491 & ~n3516 ;
  assign n3518 = n3517 ^ n3515 ;
  assign n3519 = n3518 ^ x185 ;
  assign n3521 = n3520 ^ n3519 ;
  assign n3654 = n3653 ^ n3521 ;
  assign n3655 = ~n3652 & n3654 ;
  assign n3656 = n3655 ^ n2011 ;
  assign n3839 = n3838 ^ n3656 ;
  assign n3841 = n3839 ^ x206 ;
  assign n3840 = n3839 ^ n3832 ;
  assign n3842 = n3841 ^ n3840 ;
  assign n3843 = ~n3837 & n3842 ;
  assign n3844 = n3843 ^ n3841 ;
  assign n4001 = n3844 ^ x205 ;
  assign n4002 = n4000 & n4001 ;
  assign n3657 = n3656 ^ n3651 ;
  assign n3658 = n3656 ^ n1493 ;
  assign n3659 = n3657 & n3658 ;
  assign n3660 = n3659 ^ n1493 ;
  assign n3845 = n3660 ^ n1556 ;
  assign n3661 = n2922 ^ n2050 ;
  assign n3522 = n3521 ^ n3497 ;
  assign n3523 = n3521 ^ n2900 ;
  assign n3524 = n3522 & n3523 ;
  assign n3525 = n3524 ^ n2900 ;
  assign n3662 = n3525 ^ n2922 ;
  assign n3543 = n3520 ^ n3513 ;
  assign n3544 = ~n3518 & ~n3543 ;
  assign n3541 = n3520 ^ n3518 ;
  assign n3542 = x185 & ~n3541 ;
  assign n3545 = n3544 ^ n3542 ;
  assign n3532 = n2805 ^ n2454 ;
  assign n3536 = n3509 ^ n2756 ;
  assign n3537 = n3508 & n3536 ;
  assign n3533 = n2541 ^ n2521 ;
  assign n3534 = n3533 ^ n2805 ;
  assign n3535 = n3534 ^ n3509 ;
  assign n3538 = n3537 ^ n3535 ;
  assign n3539 = ~n3532 & ~n3538 ;
  assign n3529 = n2404 ^ x184 ;
  assign n3530 = n3529 ^ n2799 ;
  assign n3526 = n3512 ^ n3501 ;
  assign n3527 = n3512 ^ n2404 ;
  assign n3528 = n3526 & ~n3527 ;
  assign n3531 = n3530 ^ n3528 ;
  assign n3540 = n3539 ^ n3531 ;
  assign n3546 = n3545 ^ n3540 ;
  assign n3663 = n3662 ^ n3546 ;
  assign n3664 = n3661 & n3663 ;
  assign n3665 = n3664 ^ n2050 ;
  assign n3846 = n3845 ^ n3665 ;
  assign n3848 = n3846 ^ x205 ;
  assign n3847 = n3846 ^ n3839 ;
  assign n3849 = n3848 ^ n3847 ;
  assign n3850 = n3844 & ~n3849 ;
  assign n3851 = n3850 ^ n3848 ;
  assign n4003 = n3851 ^ x204 ;
  assign n4004 = ~n4002 & ~n4003 ;
  assign n3666 = n3665 ^ n3660 ;
  assign n3667 = n3665 ^ n1556 ;
  assign n3668 = ~n3666 & ~n3667 ;
  assign n3669 = n3668 ^ n1556 ;
  assign n3852 = n3669 ^ n1606 ;
  assign n3670 = n2948 ^ n2091 ;
  assign n3550 = n2948 ^ n2922 ;
  assign n3547 = n3546 ^ n3525 ;
  assign n3548 = n3546 ^ n2922 ;
  assign n3549 = ~n3547 & ~n3548 ;
  assign n3551 = n3550 ^ n3549 ;
  assign n3435 = n2568 ^ x167 ;
  assign n3671 = n3551 ^ n3435 ;
  assign n3672 = n3670 & n3671 ;
  assign n3673 = n3672 ^ n2091 ;
  assign n3853 = n3852 ^ n3673 ;
  assign n3855 = n3853 ^ x204 ;
  assign n3854 = n3853 ^ n3846 ;
  assign n3856 = n3855 ^ n3854 ;
  assign n3857 = n3851 & ~n3856 ;
  assign n3858 = n3857 ^ n3855 ;
  assign n4005 = n3858 ^ x203 ;
  assign n4006 = n4004 & n4005 ;
  assign n3674 = n3673 ^ n3669 ;
  assign n3675 = n3673 ^ n1606 ;
  assign n3676 = n3674 & ~n3675 ;
  assign n3677 = n3676 ^ n1606 ;
  assign n3859 = n3677 ^ n1663 ;
  assign n3678 = n2965 ^ n2133 ;
  assign n3436 = n3435 ^ n2948 ;
  assign n3552 = n3436 & n3551 ;
  assign n3553 = n3552 ^ n2948 ;
  assign n3679 = n3553 ^ n2965 ;
  assign n3680 = n3679 ^ n2606 ;
  assign n3681 = n3678 & ~n3680 ;
  assign n3682 = n3681 ^ n2133 ;
  assign n3860 = n3859 ^ n3682 ;
  assign n3862 = n3860 ^ x203 ;
  assign n3861 = n3860 ^ n3853 ;
  assign n3863 = n3862 ^ n3861 ;
  assign n3864 = ~n3858 & n3863 ;
  assign n3865 = n3864 ^ n3862 ;
  assign n4007 = n3865 ^ x202 ;
  assign n4008 = n4006 & n4007 ;
  assign n3683 = n3682 ^ n3677 ;
  assign n3684 = n3682 ^ n1663 ;
  assign n3685 = n3683 & ~n3684 ;
  assign n3686 = n3685 ^ n1663 ;
  assign n3866 = n3686 ^ n1721 ;
  assign n3687 = n2986 ^ n2176 ;
  assign n3557 = n2648 ^ n2606 ;
  assign n3434 = n2965 ^ n2606 ;
  assign n3554 = n3553 ^ n2606 ;
  assign n3555 = ~n3434 & n3554 ;
  assign n3433 = n2986 ^ n2965 ;
  assign n3556 = n3555 ^ n3433 ;
  assign n3688 = n3557 ^ n3556 ;
  assign n3689 = ~n3687 & n3688 ;
  assign n3690 = n3689 ^ n2176 ;
  assign n3867 = n3866 ^ n3690 ;
  assign n3869 = n3867 ^ x202 ;
  assign n3868 = n3867 ^ n3860 ;
  assign n3870 = n3869 ^ n3868 ;
  assign n3871 = ~n3865 & n3870 ;
  assign n3872 = n3871 ^ n3869 ;
  assign n4009 = n3872 ^ x201 ;
  assign n4010 = ~n4008 & n4009 ;
  assign n3691 = n3690 ^ n3686 ;
  assign n3692 = n3690 ^ n1721 ;
  assign n3693 = n3691 & n3692 ;
  assign n3694 = n3693 ^ n1721 ;
  assign n3821 = n3694 ^ n1782 ;
  assign n3562 = n2691 ^ n2649 ;
  assign n3560 = n3008 ^ n2986 ;
  assign n3558 = n3557 ^ n2986 ;
  assign n3559 = ~n3556 & n3558 ;
  assign n3561 = n3560 ^ n3559 ;
  assign n3695 = n3562 ^ n3561 ;
  assign n3696 = n3008 ^ n2212 ;
  assign n3697 = n3695 & n3696 ;
  assign n3698 = n3697 ^ n2212 ;
  assign n3822 = n3821 ^ n3698 ;
  assign n3874 = n3822 ^ x201 ;
  assign n3873 = n3867 ^ n3822 ;
  assign n3875 = n3874 ^ n3873 ;
  assign n3876 = n3872 & ~n3875 ;
  assign n3877 = n3876 ^ n3874 ;
  assign n3995 = n3877 ^ x200 ;
  assign n4038 = n4010 ^ n3995 ;
  assign n4188 = n4038 ^ n3131 ;
  assign n4189 = n3125 & ~n4188 ;
  assign n4190 = n4189 ^ n3131 ;
  assign n4328 = n4190 ^ n2597 ;
  assign n4650 = n4328 ^ x231 ;
  assign n4329 = x231 & ~n4328 ;
  assign n4651 = n4329 ^ x230 ;
  assign n3432 = n2736 ^ n2692 ;
  assign n3703 = n3432 ^ n3025 ;
  assign n3563 = n3562 ^ n3008 ;
  assign n3564 = ~n3561 & ~n3563 ;
  assign n3565 = n3564 ^ n3008 ;
  assign n3704 = n3703 ^ n3565 ;
  assign n3705 = ~n3045 & n3704 ;
  assign n3706 = n3705 ^ n2254 ;
  assign n3880 = n3706 ^ n1841 ;
  assign n3699 = n3698 ^ n3694 ;
  assign n3700 = n3698 ^ n1782 ;
  assign n3701 = ~n3699 & n3700 ;
  assign n3702 = n3701 ^ n1782 ;
  assign n3881 = n3880 ^ n3702 ;
  assign n3823 = n3822 ^ x200 ;
  assign n3878 = n3823 & ~n3877 ;
  assign n3879 = n3878 ^ x200 ;
  assign n3882 = n3881 ^ n3879 ;
  assign n4012 = n3882 ^ x215 ;
  assign n4011 = n3995 & ~n4010 ;
  assign n4042 = n4012 ^ n4011 ;
  assign n4039 = n3131 ^ n3125 ;
  assign n4040 = ~n4038 & ~n4039 ;
  assign n4041 = n4040 ^ n3157 ;
  assign n4193 = n4042 ^ n4041 ;
  assign n4194 = n3169 & n4193 ;
  assign n4195 = n4194 ^ n2600 ;
  assign n4191 = n2597 & ~n4190 ;
  assign n4192 = n4191 ^ n1571 ;
  assign n4327 = n4195 ^ n4192 ;
  assign n4652 = n4651 ^ n4327 ;
  assign n4653 = ~n4650 & n4652 ;
  assign n4330 = n4329 ^ n4327 ;
  assign n4196 = n4195 ^ n4191 ;
  assign n4197 = ~n4192 & n4196 ;
  assign n4198 = n4197 ^ n1571 ;
  assign n4324 = n4198 ^ n1620 ;
  assign n4043 = n4042 ^ n4040 ;
  assign n4044 = ~n4041 & n4043 ;
  assign n4045 = n4044 ^ n3157 ;
  assign n4199 = n4045 ^ n3196 ;
  assign n4013 = n4011 & ~n4012 ;
  assign n3707 = n3706 ^ n3702 ;
  assign n3574 = n2781 ^ n2737 ;
  assign n3566 = n3565 ^ n3432 ;
  assign n3567 = n3064 ^ n3051 ;
  assign n3568 = n3567 ^ n3025 ;
  assign n3569 = n3568 ^ n3432 ;
  assign n3570 = n3569 ^ n3567 ;
  assign n3571 = n3566 & n3570 ;
  assign n3572 = n3571 ^ n3568 ;
  assign n3627 = n3574 ^ n3572 ;
  assign n3628 = ~n3051 & ~n3627 ;
  assign n3629 = n3628 ^ n3064 ;
  assign n3708 = n3629 ^ n1841 ;
  assign n3709 = n3708 ^ n3629 ;
  assign n3710 = n3709 ^ n3702 ;
  assign n3711 = ~n3707 & ~n3710 ;
  assign n3712 = n3711 ^ n3708 ;
  assign n3883 = n3712 ^ n1872 ;
  assign n3884 = n3883 ^ x215 ;
  assign n3885 = n3884 ^ n3879 ;
  assign n3886 = n3885 ^ n3883 ;
  assign n3887 = n3882 & n3886 ;
  assign n3888 = n3887 ^ n3884 ;
  assign n3994 = n3888 ^ x214 ;
  assign n4046 = n4013 ^ n3994 ;
  assign n4200 = n4199 ^ n4046 ;
  assign n4201 = n3232 & ~n4200 ;
  assign n4202 = n4201 ^ n2635 ;
  assign n4325 = n4324 ^ n4202 ;
  assign n4331 = n4325 ^ x230 ;
  assign n4332 = n4331 ^ n4325 ;
  assign n4333 = n4332 ^ n4327 ;
  assign n4334 = ~n4330 & n4333 ;
  assign n4335 = n4334 ^ n4331 ;
  assign n4654 = n4335 ^ x229 ;
  assign n4655 = n4653 & n4654 ;
  assign n4326 = n4325 ^ x229 ;
  assign n4336 = n4326 & ~n4335 ;
  assign n4337 = n4336 ^ x229 ;
  assign n4656 = n4337 ^ x228 ;
  assign n4203 = n4202 ^ n4198 ;
  assign n4204 = n4202 ^ n1620 ;
  assign n4205 = ~n4203 & ~n4204 ;
  assign n4206 = n4205 ^ n1620 ;
  assign n4322 = n4206 ^ n1676 ;
  assign n4047 = n4046 ^ n4045 ;
  assign n4014 = ~n3994 & n4013 ;
  assign n3630 = n3629 ^ n1872 ;
  assign n3713 = n3630 & ~n3712 ;
  assign n3714 = n3713 ^ n1872 ;
  assign n3889 = n3714 ^ n1916 ;
  assign n3715 = n3070 ^ n2337 ;
  assign n3573 = n2823 ^ n2782 ;
  assign n3576 = n3573 ^ n3567 ;
  assign n3575 = n3574 ^ n3573 ;
  assign n3577 = n3576 ^ n3575 ;
  assign n3578 = ~n3572 & n3577 ;
  assign n3579 = n3578 ^ n3576 ;
  assign n3716 = n3579 ^ n3070 ;
  assign n3717 = n3715 & ~n3716 ;
  assign n3718 = n3717 ^ n2337 ;
  assign n3890 = n3889 ^ n3718 ;
  assign n3892 = n3890 ^ x214 ;
  assign n3891 = n3890 ^ n3883 ;
  assign n3893 = n3892 ^ n3891 ;
  assign n3894 = n3888 & ~n3893 ;
  assign n3895 = n3894 ^ n3892 ;
  assign n3993 = n3895 ^ x213 ;
  assign n4036 = n4014 ^ n3993 ;
  assign n4048 = n4036 ^ n3196 ;
  assign n4049 = n4048 ^ n4045 ;
  assign n4050 = n4049 ^ n4036 ;
  assign n4051 = ~n4047 & n4050 ;
  assign n4052 = n4051 ^ n4048 ;
  assign n4207 = n4052 ^ n3237 ;
  assign n4208 = ~n3251 & n4207 ;
  assign n4209 = n4208 ^ n2682 ;
  assign n4323 = n4322 ^ n4209 ;
  assign n4657 = n4656 ^ n4323 ;
  assign n4658 = n4655 & n4657 ;
  assign n4338 = n4337 ^ n4323 ;
  assign n4210 = n4209 ^ n4206 ;
  assign n4211 = n4209 ^ n1676 ;
  assign n4212 = n4210 & n4211 ;
  assign n4213 = n4212 ^ n1676 ;
  assign n4339 = n4213 ^ n1733 ;
  assign n4037 = n4036 ^ n3237 ;
  assign n4053 = ~n4037 & ~n4052 ;
  assign n4054 = n4053 ^ n3237 ;
  assign n4214 = n4054 ^ n3280 ;
  assign n4015 = ~n3993 & n4014 ;
  assign n3719 = n3718 ^ n3714 ;
  assign n3720 = n3718 ^ n1916 ;
  assign n3721 = ~n3719 & n3720 ;
  assign n3722 = n3721 ^ n1916 ;
  assign n3896 = n3722 ^ n1956 ;
  assign n3585 = n2844 ^ n2824 ;
  assign n3581 = n3091 ^ n3070 ;
  assign n3580 = n3573 ^ n3091 ;
  assign n3582 = n3581 ^ n3580 ;
  assign n3583 = ~n3579 & ~n3582 ;
  assign n3584 = n3583 ^ n3581 ;
  assign n3614 = n3585 ^ n3584 ;
  assign n3723 = n3091 ^ n2379 ;
  assign n3724 = ~n3614 & n3723 ;
  assign n3725 = n3724 ^ n2379 ;
  assign n3897 = n3896 ^ n3725 ;
  assign n3899 = n3897 ^ x213 ;
  assign n3898 = n3897 ^ n3890 ;
  assign n3900 = n3899 ^ n3898 ;
  assign n3901 = n3895 & ~n3900 ;
  assign n3902 = n3901 ^ n3899 ;
  assign n3992 = n3902 ^ x212 ;
  assign n4055 = n4015 ^ n3992 ;
  assign n4215 = n4214 ^ n4055 ;
  assign n4216 = n3318 & n4215 ;
  assign n4217 = n4216 ^ n2727 ;
  assign n4340 = n4339 ^ n4217 ;
  assign n4341 = n4340 ^ x228 ;
  assign n4342 = n4341 ^ n4323 ;
  assign n4343 = n4342 ^ n4340 ;
  assign n4344 = ~n4338 & n4343 ;
  assign n4345 = n4344 ^ n4341 ;
  assign n4659 = n4345 ^ x227 ;
  assign n4660 = n4658 & n4659 ;
  assign n4218 = n4217 ^ n4213 ;
  assign n4219 = n4217 ^ n1733 ;
  assign n4220 = n4218 & ~n4219 ;
  assign n4221 = n4220 ^ n1733 ;
  assign n4346 = n4221 ^ n1795 ;
  assign n4056 = n4055 ^ n4054 ;
  assign n4057 = n4055 ^ n3280 ;
  assign n4058 = ~n4056 & n4057 ;
  assign n4059 = n4058 ^ n3280 ;
  assign n4222 = n4059 ^ n3323 ;
  assign n4016 = n3992 & n4015 ;
  assign n3726 = n3725 ^ n3722 ;
  assign n3727 = n3725 ^ n1956 ;
  assign n3728 = ~n3726 & ~n3727 ;
  assign n3729 = n3728 ^ n1956 ;
  assign n3903 = n3729 ^ n1997 ;
  assign n3730 = n3111 ^ n2424 ;
  assign n3592 = n2865 ^ n2845 ;
  assign n3587 = n3111 ^ n3091 ;
  assign n3586 = n3585 ^ n3111 ;
  assign n3588 = n3587 ^ n3586 ;
  assign n3589 = n3584 & n3588 ;
  assign n3590 = n3589 ^ n3587 ;
  assign n3731 = n3592 ^ n3590 ;
  assign n3732 = n3730 & ~n3731 ;
  assign n3733 = n3732 ^ n2424 ;
  assign n3904 = n3903 ^ n3733 ;
  assign n3906 = n3904 ^ x212 ;
  assign n3905 = n3904 ^ n3897 ;
  assign n3907 = n3906 ^ n3905 ;
  assign n3908 = ~n3902 & n3907 ;
  assign n3909 = n3908 ^ n3906 ;
  assign n3991 = n3909 ^ x211 ;
  assign n4060 = n4016 ^ n3991 ;
  assign n4223 = n4222 ^ n4060 ;
  assign n4224 = ~n3337 & n4223 ;
  assign n4225 = n4224 ^ n2772 ;
  assign n4347 = n4346 ^ n4225 ;
  assign n4349 = n4347 ^ x227 ;
  assign n4348 = n4347 ^ n4340 ;
  assign n4350 = n4349 ^ n4348 ;
  assign n4351 = ~n4345 & n4350 ;
  assign n4352 = n4351 ^ n4349 ;
  assign n4661 = n4352 ^ x226 ;
  assign n4662 = n4660 & ~n4661 ;
  assign n4226 = n4225 ^ n4221 ;
  assign n4227 = n4225 ^ n1795 ;
  assign n4228 = n4226 & n4227 ;
  assign n4229 = n4228 ^ n1795 ;
  assign n4353 = n4229 ^ n1853 ;
  assign n4061 = n4060 ^ n4059 ;
  assign n4017 = ~n3991 & ~n4016 ;
  assign n3734 = n3733 ^ n3729 ;
  assign n3735 = n3733 ^ n1997 ;
  assign n3736 = ~n3734 & n3735 ;
  assign n3737 = n3736 ^ n1997 ;
  assign n3910 = n3737 ^ n2043 ;
  assign n3738 = n3145 ^ n2464 ;
  assign n3591 = n2887 ^ n2866 ;
  assign n3594 = n3591 ^ n3111 ;
  assign n3593 = n3592 ^ n3591 ;
  assign n3595 = n3594 ^ n3593 ;
  assign n3596 = ~n3590 & n3595 ;
  assign n3597 = n3596 ^ n3594 ;
  assign n3739 = n3597 ^ n3145 ;
  assign n3740 = ~n3738 & ~n3739 ;
  assign n3741 = n3740 ^ n2464 ;
  assign n3911 = n3910 ^ n3741 ;
  assign n3913 = n3911 ^ x211 ;
  assign n3912 = n3911 ^ n3904 ;
  assign n3914 = n3913 ^ n3912 ;
  assign n3915 = ~n3909 & n3914 ;
  assign n3916 = n3915 ^ n3913 ;
  assign n3990 = n3916 ^ x210 ;
  assign n4034 = n4017 ^ n3990 ;
  assign n4062 = n4034 ^ n3323 ;
  assign n4063 = n4062 ^ n4034 ;
  assign n4064 = n4063 ^ n4059 ;
  assign n4065 = n4061 & ~n4064 ;
  assign n4066 = n4065 ^ n4062 ;
  assign n4230 = n4066 ^ n3363 ;
  assign n4231 = n3401 & ~n4230 ;
  assign n4232 = n4231 ^ n2814 ;
  assign n4354 = n4353 ^ n4232 ;
  assign n4356 = n4354 ^ x226 ;
  assign n4355 = n4354 ^ n4347 ;
  assign n4357 = n4356 ^ n4355 ;
  assign n4358 = n4352 & ~n4357 ;
  assign n4359 = n4358 ^ n4356 ;
  assign n4663 = n4359 ^ x225 ;
  assign n4664 = n4662 & ~n4663 ;
  assign n4233 = n4232 ^ n4229 ;
  assign n4234 = n4232 ^ n1853 ;
  assign n4235 = n4233 & ~n4234 ;
  assign n4236 = n4235 ^ n1853 ;
  assign n4360 = n4236 ^ n2833 ;
  assign n4035 = n4034 ^ n3363 ;
  assign n4067 = n4035 & ~n4066 ;
  assign n4068 = n4067 ^ n3363 ;
  assign n4237 = n4068 ^ n3406 ;
  assign n4018 = n3990 & n4017 ;
  assign n3742 = n3741 ^ n3737 ;
  assign n3743 = n3741 ^ n2043 ;
  assign n3744 = n3742 & ~n3743 ;
  assign n3745 = n3744 ^ n2043 ;
  assign n3917 = n3745 ^ n2083 ;
  assign n3746 = n3181 ^ n2484 ;
  assign n3603 = n2909 ^ n2888 ;
  assign n3599 = n3181 ^ n3145 ;
  assign n3598 = n3591 ^ n3181 ;
  assign n3600 = n3599 ^ n3598 ;
  assign n3601 = n3597 & ~n3600 ;
  assign n3602 = n3601 ^ n3599 ;
  assign n3747 = n3603 ^ n3602 ;
  assign n3748 = n3746 & ~n3747 ;
  assign n3749 = n3748 ^ n2484 ;
  assign n3918 = n3917 ^ n3749 ;
  assign n3920 = n3918 ^ x210 ;
  assign n3919 = n3918 ^ n3911 ;
  assign n3921 = n3920 ^ n3919 ;
  assign n3922 = n3916 & ~n3921 ;
  assign n3923 = n3922 ^ n3920 ;
  assign n3989 = n3923 ^ x209 ;
  assign n4069 = n4018 ^ n3989 ;
  assign n4238 = n4237 ^ n4069 ;
  assign n4239 = ~n3437 & ~n4238 ;
  assign n4240 = n4239 ^ n2835 ;
  assign n4361 = n4360 ^ n4240 ;
  assign n4363 = n4361 ^ x225 ;
  assign n4362 = n4361 ^ n4354 ;
  assign n4364 = n4363 ^ n4362 ;
  assign n4365 = n4359 & ~n4364 ;
  assign n4366 = n4365 ^ n4363 ;
  assign n4665 = n4366 ^ x224 ;
  assign n4666 = n4664 & n4665 ;
  assign n4241 = n4240 ^ n4236 ;
  assign n4242 = n4240 ^ n2833 ;
  assign n4243 = n4241 & n4242 ;
  assign n4244 = n4243 ^ n2833 ;
  assign n4367 = n4244 ^ n1929 ;
  assign n4070 = n4069 ^ n4068 ;
  assign n4071 = n4069 ^ n3406 ;
  assign n4072 = n4070 & n4071 ;
  assign n4073 = n4072 ^ n3406 ;
  assign n4245 = n4073 ^ n3637 ;
  assign n4019 = ~n3989 & ~n4018 ;
  assign n3750 = n3749 ^ n3745 ;
  assign n3751 = n3749 ^ n2083 ;
  assign n3752 = ~n3750 & ~n3751 ;
  assign n3753 = n3752 ^ n2083 ;
  assign n3924 = n3753 ^ n2120 ;
  assign n3609 = n2931 ^ n2910 ;
  assign n3605 = n3217 ^ n3181 ;
  assign n3604 = n3603 ^ n3217 ;
  assign n3606 = n3605 ^ n3604 ;
  assign n3607 = n3602 & ~n3606 ;
  assign n3608 = n3607 ^ n3605 ;
  assign n3610 = n3609 ^ n3608 ;
  assign n3754 = n3216 & n3610 ;
  assign n3755 = n3754 ^ n2505 ;
  assign n3925 = n3924 ^ n3755 ;
  assign n3927 = n3925 ^ x209 ;
  assign n3926 = n3925 ^ n3918 ;
  assign n3928 = n3927 ^ n3926 ;
  assign n3929 = n3923 & ~n3928 ;
  assign n3930 = n3929 ^ n3927 ;
  assign n3988 = n3930 ^ x208 ;
  assign n4032 = n4019 ^ n3988 ;
  assign n4246 = n4245 ^ n4032 ;
  assign n4247 = n3466 & ~n4246 ;
  assign n4248 = n4247 ^ n2856 ;
  assign n4368 = n4367 ^ n4248 ;
  assign n4370 = n4368 ^ x224 ;
  assign n4369 = n4368 ^ n4361 ;
  assign n4371 = n4370 ^ n4369 ;
  assign n4372 = ~n4366 & n4371 ;
  assign n4373 = n4372 ^ n4370 ;
  assign n4667 = n4373 ^ x239 ;
  assign n4668 = ~n4666 & n4667 ;
  assign n4249 = n4248 ^ n4244 ;
  assign n4250 = n4248 ^ n1929 ;
  assign n4251 = ~n4249 & n4250 ;
  assign n4252 = n4251 ^ n1929 ;
  assign n4374 = n4252 ^ n1970 ;
  assign n4033 = n4032 ^ n3637 ;
  assign n4074 = n4073 ^ n4032 ;
  assign n4075 = ~n4033 & ~n4074 ;
  assign n4076 = n4075 ^ n3637 ;
  assign n4253 = n4076 ^ n3645 ;
  assign n4020 = n3988 & n4019 ;
  assign n3756 = n3755 ^ n3753 ;
  assign n3622 = n2952 ^ n2932 ;
  assign n3616 = n3263 ^ n2527 ;
  assign n3618 = n3616 ^ n3217 ;
  assign n3617 = n3616 ^ n3609 ;
  assign n3619 = n3618 ^ n3617 ;
  assign n3620 = ~n3608 & n3619 ;
  assign n3621 = n3620 ^ n3618 ;
  assign n3623 = n3622 ^ n3621 ;
  assign n3624 = n3263 & ~n3623 ;
  assign n3625 = n3624 ^ n2527 ;
  assign n3757 = n3625 ^ n2120 ;
  assign n3758 = n3757 ^ n3625 ;
  assign n3759 = n3758 ^ n3753 ;
  assign n3760 = ~n3756 & ~n3759 ;
  assign n3761 = n3760 ^ n3757 ;
  assign n3931 = n3761 ^ n2163 ;
  assign n3933 = n3931 ^ x208 ;
  assign n3932 = n3931 ^ n3925 ;
  assign n3934 = n3933 ^ n3932 ;
  assign n3935 = ~n3930 & n3934 ;
  assign n3936 = n3935 ^ n3933 ;
  assign n3987 = n3936 ^ x223 ;
  assign n4077 = n4020 ^ n3987 ;
  assign n4254 = n4253 ^ n4077 ;
  assign n4255 = n3495 & n4254 ;
  assign n4256 = n4255 ^ n2878 ;
  assign n4375 = n4374 ^ n4256 ;
  assign n4377 = n4375 ^ x239 ;
  assign n4376 = n4375 ^ n4368 ;
  assign n4378 = n4377 ^ n4376 ;
  assign n4379 = n4373 & ~n4378 ;
  assign n4380 = n4379 ^ n4377 ;
  assign n4669 = n4380 ^ x238 ;
  assign n4670 = ~n4668 & n4669 ;
  assign n4257 = n4256 ^ n4252 ;
  assign n4258 = n4256 ^ n1970 ;
  assign n4259 = n4257 & ~n4258 ;
  assign n4260 = n4259 ^ n1970 ;
  assign n4381 = n4260 ^ n2011 ;
  assign n4078 = n4077 ^ n4076 ;
  assign n4079 = n4077 ^ n3645 ;
  assign n4080 = ~n4078 & ~n4079 ;
  assign n4081 = n4080 ^ n3645 ;
  assign n4261 = n4081 ^ n3654 ;
  assign n4021 = ~n3987 & n4020 ;
  assign n3626 = n3625 ^ n2163 ;
  assign n3762 = ~n3626 & n3761 ;
  assign n3763 = n3762 ^ n2163 ;
  assign n3937 = n3763 ^ n2571 ;
  assign n3764 = n3302 ^ n3295 ;
  assign n3765 = n2974 ^ n2953 ;
  assign n3767 = n3765 ^ n3616 ;
  assign n3766 = n3765 ^ n3622 ;
  assign n3768 = n3767 ^ n3766 ;
  assign n3769 = n3621 & n3768 ;
  assign n3770 = n3769 ^ n3767 ;
  assign n3771 = n3770 ^ n3302 ;
  assign n3772 = n3764 & n3771 ;
  assign n3773 = n3772 ^ n3295 ;
  assign n3938 = n3937 ^ n3773 ;
  assign n3940 = n3938 ^ x223 ;
  assign n3939 = n3938 ^ n3931 ;
  assign n3941 = n3940 ^ n3939 ;
  assign n3942 = n3936 & ~n3941 ;
  assign n3943 = n3942 ^ n3940 ;
  assign n3986 = n3943 ^ x222 ;
  assign n4030 = n4021 ^ n3986 ;
  assign n4262 = n4261 ^ n4030 ;
  assign n4263 = ~n3522 & ~n4262 ;
  assign n4264 = n4263 ^ n2900 ;
  assign n4382 = n4381 ^ n4264 ;
  assign n4384 = n4382 ^ x238 ;
  assign n4383 = n4382 ^ n4375 ;
  assign n4385 = n4384 ^ n4383 ;
  assign n4386 = ~n4380 & n4385 ;
  assign n4387 = n4386 ^ n4384 ;
  assign n4649 = n4387 ^ x237 ;
  assign n4722 = n4670 ^ n4649 ;
  assign n3431 = n3428 ^ n3427 ;
  assign n3611 = n3610 ^ n3431 ;
  assign n3613 = n3420 ^ n3419 ;
  assign n3615 = n3614 ^ n3613 ;
  assign n4144 = n2411 ^ x216 ;
  assign n4145 = n4144 ^ n3532 ;
  assign n3807 = n3455 ^ n2665 ;
  assign n3813 = n3039 ^ n3018 ;
  assign n3780 = n3352 ^ n3302 ;
  assign n3779 = n3765 ^ n3352 ;
  assign n3781 = n3780 ^ n3779 ;
  assign n3782 = n3770 & ~n3781 ;
  assign n3783 = n3782 ^ n3780 ;
  assign n3794 = n3391 ^ n3352 ;
  assign n3784 = n2995 ^ n2975 ;
  assign n3793 = n3784 ^ n3391 ;
  assign n3795 = n3794 ^ n3793 ;
  assign n3796 = ~n3783 & n3795 ;
  assign n3797 = n3796 ^ n3794 ;
  assign n3809 = n3455 ^ n3391 ;
  assign n3798 = n3017 ^ n2996 ;
  assign n3808 = n3798 ^ n3455 ;
  assign n3810 = n3809 ^ n3808 ;
  assign n3811 = ~n3797 & ~n3810 ;
  assign n3812 = n3811 ^ n3809 ;
  assign n3814 = n3813 ^ n3812 ;
  assign n3815 = n3807 & ~n3814 ;
  assign n3816 = n3815 ^ n2665 ;
  assign n3792 = n3391 ^ n2618 ;
  assign n3799 = n3798 ^ n3797 ;
  assign n3800 = ~n3792 & ~n3799 ;
  assign n3801 = n3800 ^ n2618 ;
  assign n3778 = n3352 ^ n2580 ;
  assign n3785 = n3784 ^ n3783 ;
  assign n3786 = n3778 & ~n3785 ;
  assign n3787 = n3786 ^ n2580 ;
  assign n3774 = n3773 ^ n3763 ;
  assign n3775 = n3773 ^ n2571 ;
  assign n3776 = n3774 & ~n3775 ;
  assign n3777 = n3776 ^ n2571 ;
  assign n3788 = n3787 ^ n3777 ;
  assign n3789 = n3787 ^ n2573 ;
  assign n3790 = ~n3788 & ~n3789 ;
  assign n3791 = n3790 ^ n2573 ;
  assign n3802 = n3801 ^ n3791 ;
  assign n3803 = n3801 ^ n2283 ;
  assign n3804 = n3802 & ~n3803 ;
  assign n3805 = n3804 ^ n2283 ;
  assign n3959 = n3816 ^ n3805 ;
  assign n3960 = n3483 ^ n2710 ;
  assign n3966 = n3061 ^ n3040 ;
  assign n3962 = n3483 ^ n3455 ;
  assign n3961 = n3813 ^ n3483 ;
  assign n3963 = n3962 ^ n3961 ;
  assign n3964 = ~n3812 & n3963 ;
  assign n3965 = n3964 ^ n3962 ;
  assign n3967 = n3966 ^ n3965 ;
  assign n3968 = n3960 & n3967 ;
  assign n3969 = n3968 ^ n2710 ;
  assign n3970 = n3969 ^ n2325 ;
  assign n3971 = n3970 ^ n3969 ;
  assign n3972 = n3971 ^ n3805 ;
  assign n3973 = n3959 & ~n3972 ;
  assign n3974 = n3973 ^ n3970 ;
  assign n4105 = n3510 ^ n2756 ;
  assign n4111 = n3084 ^ n3062 ;
  assign n4107 = n3510 ^ n3483 ;
  assign n4106 = n3966 ^ n3510 ;
  assign n4108 = n4107 ^ n4106 ;
  assign n4109 = ~n3965 & n4108 ;
  assign n4110 = n4109 ^ n4107 ;
  assign n4112 = n4111 ^ n4110 ;
  assign n4113 = ~n4105 & n4112 ;
  assign n4114 = n4113 ^ n2756 ;
  assign n4116 = n4114 ^ n2362 ;
  assign n4115 = n4114 ^ n3969 ;
  assign n4117 = n4116 ^ n4115 ;
  assign n4118 = n3974 & ~n4117 ;
  assign n4119 = n4118 ^ n4116 ;
  assign n4142 = n4114 ^ n2411 ;
  assign n4143 = ~n4119 & n4142 ;
  assign n4146 = n4145 ^ n4143 ;
  assign n4134 = n3538 ^ n2805 ;
  assign n4138 = n4111 ^ n3510 ;
  assign n4139 = ~n4110 & ~n4138 ;
  assign n4135 = n3538 ^ n3085 ;
  assign n4136 = n4135 ^ n3104 ;
  assign n4137 = n4136 ^ n4111 ;
  assign n4140 = n4139 ^ n4137 ;
  assign n4141 = n4134 & ~n4140 ;
  assign n4147 = n4146 ^ n4141 ;
  assign n3818 = n3791 ^ n2283 ;
  assign n3819 = n3818 ^ n3801 ;
  assign n3820 = n3819 ^ x220 ;
  assign n3944 = n3777 ^ n2573 ;
  assign n3945 = n3944 ^ n3787 ;
  assign n3947 = n3945 ^ x222 ;
  assign n3946 = n3945 ^ n3938 ;
  assign n3948 = n3947 ^ n3946 ;
  assign n3949 = n3943 & ~n3948 ;
  assign n3950 = n3949 ^ n3947 ;
  assign n3952 = n3819 ^ x221 ;
  assign n3951 = n3945 ^ n3819 ;
  assign n3953 = n3952 ^ n3951 ;
  assign n3954 = n3950 & ~n3953 ;
  assign n3955 = n3954 ^ n3952 ;
  assign n3956 = n3820 & ~n3955 ;
  assign n3957 = n3956 ^ x220 ;
  assign n3806 = n3805 ^ n2325 ;
  assign n3817 = n3816 ^ n3806 ;
  assign n3958 = n3957 ^ n3817 ;
  assign n3975 = n3974 ^ n2362 ;
  assign n3976 = n3975 ^ x219 ;
  assign n3977 = n3976 ^ n3817 ;
  assign n3978 = n3977 ^ n3975 ;
  assign n3979 = n3958 & ~n3978 ;
  assign n3980 = n3979 ^ n3976 ;
  assign n3981 = n3980 ^ x218 ;
  assign n3982 = n3957 ^ x219 ;
  assign n3983 = n3982 ^ n3817 ;
  assign n3984 = n3955 ^ x220 ;
  assign n3985 = n3950 ^ x221 ;
  assign n4022 = ~n3986 & n4021 ;
  assign n4023 = ~n3985 & n4022 ;
  assign n4024 = ~n3984 & ~n4023 ;
  assign n4025 = ~n3983 & ~n4024 ;
  assign n4122 = n3981 & ~n4025 ;
  assign n4120 = n4119 ^ n2411 ;
  assign n4128 = n4122 ^ n4120 ;
  assign n4101 = n3975 ^ x218 ;
  assign n4102 = n3980 & ~n4101 ;
  assign n4103 = n4102 ^ x218 ;
  assign n4131 = n4120 ^ n4103 ;
  assign n4132 = n4128 & ~n4131 ;
  assign n4129 = n4128 ^ n4103 ;
  assign n4130 = ~x217 & ~n4129 ;
  assign n4133 = n4132 ^ n4130 ;
  assign n4148 = n4147 ^ n4133 ;
  assign n4104 = n4103 ^ x217 ;
  assign n4121 = n4120 ^ n4104 ;
  assign n4123 = n4122 ^ n4121 ;
  assign n4026 = n4025 ^ n3981 ;
  assign n4027 = n4026 ^ n3688 ;
  assign n4093 = n4024 ^ n3983 ;
  assign n4028 = n4023 ^ n3984 ;
  assign n4029 = n4028 ^ n3671 ;
  assign n4085 = n4022 ^ n3985 ;
  assign n4031 = n4030 ^ n3654 ;
  assign n4082 = n4081 ^ n4030 ;
  assign n4083 = ~n4031 & n4082 ;
  assign n4084 = n4083 ^ n3654 ;
  assign n4086 = n4085 ^ n4084 ;
  assign n4087 = n4085 ^ n3663 ;
  assign n4088 = n4086 & ~n4087 ;
  assign n4089 = n4088 ^ n3663 ;
  assign n4090 = n4089 ^ n4028 ;
  assign n4091 = ~n4029 & n4090 ;
  assign n4092 = n4091 ^ n3671 ;
  assign n4094 = n4093 ^ n4092 ;
  assign n4095 = n4093 ^ n3680 ;
  assign n4096 = ~n4094 & ~n4095 ;
  assign n4097 = n4096 ^ n3680 ;
  assign n4098 = n4097 ^ n4026 ;
  assign n4099 = n4027 & n4098 ;
  assign n4100 = n4099 ^ n3688 ;
  assign n4124 = n4123 ^ n4100 ;
  assign n4125 = n4123 ^ n3695 ;
  assign n4126 = n4124 & ~n4125 ;
  assign n4127 = n4126 ^ n3695 ;
  assign n4149 = n4148 ^ n4127 ;
  assign n4150 = n4148 ^ n3704 ;
  assign n4151 = n4149 & ~n4150 ;
  assign n4152 = n4151 ^ n3704 ;
  assign n4153 = n4152 ^ n3627 ;
  assign n4154 = n3716 ^ n3416 ;
  assign n4155 = n4154 ^ n3716 ;
  assign n4156 = n4155 ^ n4152 ;
  assign n4157 = n4153 & n4156 ;
  assign n4158 = n4157 ^ n4154 ;
  assign n4161 = n3716 ^ n3614 ;
  assign n4159 = n3418 ^ n3416 ;
  assign n4160 = n4159 ^ n3614 ;
  assign n4162 = n4161 ^ n4160 ;
  assign n4163 = ~n4158 & ~n4162 ;
  assign n4164 = n4163 ^ n4161 ;
  assign n4165 = ~n3615 & n4164 ;
  assign n4166 = n4165 ^ n3614 ;
  assign n3612 = n3422 ^ n3421 ;
  assign n4167 = n4166 ^ n3612 ;
  assign n4169 = n3739 ^ n3731 ;
  assign n4168 = n4166 ^ n3739 ;
  assign n4170 = n4169 ^ n4168 ;
  assign n4171 = n4167 & n4170 ;
  assign n4172 = n4171 ^ n4169 ;
  assign n4175 = n3747 ^ n3739 ;
  assign n4173 = n3424 ^ n3423 ;
  assign n4174 = n4173 ^ n3747 ;
  assign n4176 = n4175 ^ n4174 ;
  assign n4177 = n4172 & n4176 ;
  assign n4178 = n4177 ^ n4175 ;
  assign n4181 = n3747 ^ n3610 ;
  assign n4179 = n3426 ^ n3425 ;
  assign n4180 = n4179 ^ n3610 ;
  assign n4182 = n4181 ^ n4180 ;
  assign n4183 = n4178 & n4182 ;
  assign n4184 = n4183 ^ n4181 ;
  assign n4185 = n3611 & ~n4184 ;
  assign n4186 = n4185 ^ n3610 ;
  assign n3430 = n3429 ^ n3415 ;
  assign n4187 = n4186 ^ n3430 ;
  assign n4872 = n4654 ^ n4653 ;
  assign n4265 = n4264 ^ n4260 ;
  assign n4266 = n4264 ^ n2011 ;
  assign n4267 = ~n4265 & ~n4266 ;
  assign n4268 = n4267 ^ n2011 ;
  assign n4388 = n4268 ^ n2050 ;
  assign n4269 = n4084 ^ n3663 ;
  assign n4270 = n4269 ^ n4085 ;
  assign n4271 = n3547 & ~n4270 ;
  assign n4272 = n4271 ^ n2922 ;
  assign n4389 = n4388 ^ n4272 ;
  assign n4391 = n4389 ^ x237 ;
  assign n4390 = n4389 ^ n4382 ;
  assign n4392 = n4391 ^ n4390 ;
  assign n4393 = ~n4387 & n4392 ;
  assign n4394 = n4393 ^ n4391 ;
  assign n4273 = n4272 ^ n4268 ;
  assign n4274 = n4272 ^ n2050 ;
  assign n4275 = ~n4273 & n4274 ;
  assign n4276 = n4275 ^ n2050 ;
  assign n4395 = n4276 ^ n2091 ;
  assign n4277 = n3671 ^ n2948 ;
  assign n4278 = n4089 ^ n3671 ;
  assign n4279 = n4278 ^ n4028 ;
  assign n4280 = n4277 & ~n4279 ;
  assign n4281 = n4280 ^ n2948 ;
  assign n4396 = n4395 ^ n4281 ;
  assign n4398 = n4396 ^ x236 ;
  assign n4397 = n4396 ^ n4389 ;
  assign n4399 = n4398 ^ n4397 ;
  assign n4400 = ~n4394 & n4399 ;
  assign n4401 = n4400 ^ n4398 ;
  assign n4647 = n4401 ^ x235 ;
  assign n4648 = n4394 ^ x236 ;
  assign n4671 = ~n4649 & ~n4670 ;
  assign n4672 = n4648 & ~n4671 ;
  assign n4673 = ~n4647 & ~n4672 ;
  assign n4282 = n4281 ^ n4276 ;
  assign n4283 = n4281 ^ n2091 ;
  assign n4284 = ~n4282 & n4283 ;
  assign n4285 = n4284 ^ n2091 ;
  assign n4402 = n4285 ^ n2133 ;
  assign n4286 = n4092 ^ n3680 ;
  assign n4287 = n4286 ^ n4093 ;
  assign n4288 = ~n3554 & ~n4287 ;
  assign n4289 = n4288 ^ n2965 ;
  assign n4403 = n4402 ^ n4289 ;
  assign n4405 = n4403 ^ x235 ;
  assign n4404 = n4403 ^ n4396 ;
  assign n4406 = n4405 ^ n4404 ;
  assign n4407 = ~n4401 & n4406 ;
  assign n4408 = n4407 ^ n4405 ;
  assign n4674 = n4408 ^ x234 ;
  assign n4675 = ~n4673 & n4674 ;
  assign n4290 = n4289 ^ n4285 ;
  assign n4291 = n4289 ^ n2133 ;
  assign n4292 = ~n4290 & n4291 ;
  assign n4293 = n4292 ^ n2133 ;
  assign n4409 = n4293 ^ n2176 ;
  assign n4294 = n3688 ^ n2986 ;
  assign n4295 = n4097 ^ n3688 ;
  assign n4296 = n4295 ^ n4026 ;
  assign n4297 = ~n4294 & ~n4296 ;
  assign n4298 = n4297 ^ n2986 ;
  assign n4410 = n4409 ^ n4298 ;
  assign n4412 = n4410 ^ x234 ;
  assign n4411 = n4410 ^ n4403 ;
  assign n4413 = n4412 ^ n4411 ;
  assign n4414 = ~n4408 & n4413 ;
  assign n4415 = n4414 ^ n4412 ;
  assign n4676 = n4415 ^ x233 ;
  assign n4677 = n4675 & ~n4676 ;
  assign n4299 = n4298 ^ n4293 ;
  assign n4300 = n4298 ^ n2176 ;
  assign n4301 = n4299 & ~n4300 ;
  assign n4302 = n4301 ^ n2176 ;
  assign n4319 = n4302 ^ n2212 ;
  assign n4303 = n3695 ^ n3008 ;
  assign n4304 = n4100 ^ n3695 ;
  assign n4305 = n4304 ^ n4123 ;
  assign n4306 = n4303 & ~n4305 ;
  assign n4307 = n4306 ^ n3008 ;
  assign n4320 = n4319 ^ n4307 ;
  assign n4417 = n4320 ^ x233 ;
  assign n4416 = n4410 ^ n4320 ;
  assign n4418 = n4417 ^ n4416 ;
  assign n4419 = n4415 & ~n4418 ;
  assign n4420 = n4419 ^ n4417 ;
  assign n4678 = n4420 ^ x232 ;
  assign n4679 = ~n4677 & ~n4678 ;
  assign n4321 = n4320 ^ x232 ;
  assign n4421 = n4321 & ~n4420 ;
  assign n4422 = n4421 ^ x232 ;
  assign n4680 = n4422 ^ x247 ;
  assign n4308 = n4307 ^ n4302 ;
  assign n4309 = n4127 ^ n3704 ;
  assign n4310 = n4309 ^ n4148 ;
  assign n4311 = ~n3566 & ~n4310 ;
  assign n4312 = n4311 ^ n3025 ;
  assign n4313 = n4312 ^ n2212 ;
  assign n4314 = n4313 ^ n4312 ;
  assign n4315 = n4314 ^ n4302 ;
  assign n4316 = ~n4308 & n4315 ;
  assign n4317 = n4316 ^ n4313 ;
  assign n4318 = n4317 ^ n2254 ;
  assign n4681 = n4680 ^ n4318 ;
  assign n4682 = ~n4679 & ~n4681 ;
  assign n4423 = n4422 ^ n4318 ;
  assign n4428 = n3627 ^ n3567 ;
  assign n4429 = n3627 ^ n3416 ;
  assign n4430 = n4429 ^ n4152 ;
  assign n4431 = ~n4428 & ~n4430 ;
  assign n4432 = n4431 ^ n3567 ;
  assign n4424 = n4312 ^ n2254 ;
  assign n4425 = n4317 & ~n4424 ;
  assign n4426 = n4425 ^ n2254 ;
  assign n4427 = n4426 ^ n3064 ;
  assign n4433 = n4432 ^ n4427 ;
  assign n4434 = n4433 ^ x247 ;
  assign n4435 = n4434 ^ n4318 ;
  assign n4436 = n4435 ^ n4433 ;
  assign n4437 = n4423 & ~n4436 ;
  assign n4438 = n4437 ^ n4434 ;
  assign n4683 = n4438 ^ x246 ;
  assign n4684 = ~n4682 & n4683 ;
  assign n4444 = n4159 ^ n4158 ;
  assign n4445 = n3579 & ~n4444 ;
  assign n4446 = n4445 ^ n3070 ;
  assign n4439 = n4432 ^ n4426 ;
  assign n4440 = n4432 ^ n3064 ;
  assign n4441 = ~n4439 & ~n4440 ;
  assign n4442 = n4441 ^ n3064 ;
  assign n4443 = n4442 ^ n2337 ;
  assign n4447 = n4446 ^ n4443 ;
  assign n4449 = n4447 ^ x246 ;
  assign n4448 = n4447 ^ n4433 ;
  assign n4450 = n4449 ^ n4448 ;
  assign n4451 = n4438 & ~n4450 ;
  assign n4452 = n4451 ^ n4449 ;
  assign n4685 = n4452 ^ x245 ;
  assign n4686 = n4684 & n4685 ;
  assign n4458 = n3614 ^ n3091 ;
  assign n4459 = n4164 ^ n3613 ;
  assign n4460 = n4458 & n4459 ;
  assign n4461 = n4460 ^ n3091 ;
  assign n4453 = n4446 ^ n4442 ;
  assign n4454 = n4446 ^ n2337 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4456 = n4455 ^ n2337 ;
  assign n4457 = n4456 ^ n2379 ;
  assign n4462 = n4461 ^ n4457 ;
  assign n4464 = n4462 ^ x245 ;
  assign n4463 = n4462 ^ n4447 ;
  assign n4465 = n4464 ^ n4463 ;
  assign n4466 = n4452 & ~n4465 ;
  assign n4467 = n4466 ^ n4464 ;
  assign n4687 = n4467 ^ x244 ;
  assign n4688 = ~n4686 & ~n4687 ;
  assign n4473 = n3731 ^ n3111 ;
  assign n4474 = n4167 ^ n3731 ;
  assign n4475 = ~n4473 & n4474 ;
  assign n4476 = n4475 ^ n3111 ;
  assign n4468 = n4461 ^ n4456 ;
  assign n4469 = n4461 ^ n2379 ;
  assign n4470 = ~n4468 & n4469 ;
  assign n4471 = n4470 ^ n2379 ;
  assign n4472 = n4471 ^ n2424 ;
  assign n4477 = n4476 ^ n4472 ;
  assign n4479 = n4477 ^ x244 ;
  assign n4478 = n4477 ^ n4462 ;
  assign n4480 = n4479 ^ n4478 ;
  assign n4481 = n4467 & ~n4480 ;
  assign n4482 = n4481 ^ n4479 ;
  assign n4689 = n4482 ^ x243 ;
  assign n4690 = n4688 & ~n4689 ;
  assign n4488 = n4173 ^ n4172 ;
  assign n4489 = ~n3597 & ~n4488 ;
  assign n4490 = n4489 ^ n3145 ;
  assign n4483 = n4476 ^ n4471 ;
  assign n4484 = n4476 ^ n2424 ;
  assign n4485 = n4483 & n4484 ;
  assign n4486 = n4485 ^ n2424 ;
  assign n4487 = n4486 ^ n2464 ;
  assign n4491 = n4490 ^ n4487 ;
  assign n4493 = n4491 ^ x243 ;
  assign n4492 = n4491 ^ n4477 ;
  assign n4494 = n4493 ^ n4492 ;
  assign n4495 = n4482 & ~n4494 ;
  assign n4496 = n4495 ^ n4493 ;
  assign n4691 = n4496 ^ x242 ;
  assign n4692 = n4690 & ~n4691 ;
  assign n4502 = n3747 ^ n3181 ;
  assign n4503 = n4179 ^ n4178 ;
  assign n4504 = ~n4502 & ~n4503 ;
  assign n4505 = n4504 ^ n3181 ;
  assign n4497 = n4490 ^ n4486 ;
  assign n4498 = n4490 ^ n2464 ;
  assign n4499 = ~n4497 & ~n4498 ;
  assign n4500 = n4499 ^ n2464 ;
  assign n4501 = n4500 ^ n2484 ;
  assign n4506 = n4505 ^ n4501 ;
  assign n4508 = n4506 ^ x242 ;
  assign n4507 = n4506 ^ n4491 ;
  assign n4509 = n4508 ^ n4507 ;
  assign n4510 = n4496 & ~n4509 ;
  assign n4511 = n4510 ^ n4508 ;
  assign n4693 = n4511 ^ x241 ;
  assign n4694 = ~n4692 & n4693 ;
  assign n4517 = n4184 ^ n3431 ;
  assign n4518 = n3610 ^ n3217 ;
  assign n4519 = ~n4517 & ~n4518 ;
  assign n4520 = n4519 ^ n3217 ;
  assign n4512 = n4505 ^ n4500 ;
  assign n4513 = n4505 ^ n2484 ;
  assign n4514 = n4512 & n4513 ;
  assign n4515 = n4514 ^ n2484 ;
  assign n4516 = n4515 ^ n2505 ;
  assign n4521 = n4520 ^ n4516 ;
  assign n4523 = n4521 ^ x241 ;
  assign n4522 = n4521 ^ n4506 ;
  assign n4524 = n4523 ^ n4522 ;
  assign n4525 = n4511 & ~n4524 ;
  assign n4526 = n4525 ^ n4523 ;
  assign n4695 = n4526 ^ x240 ;
  assign n4696 = ~n4694 & n4695 ;
  assign n4527 = n4520 ^ n4515 ;
  assign n4528 = n3623 ^ n3616 ;
  assign n4529 = n3623 ^ n3430 ;
  assign n4530 = n4529 ^ n4186 ;
  assign n4531 = n4528 & ~n4530 ;
  assign n4532 = n4531 ^ n3616 ;
  assign n4533 = n4532 ^ n2505 ;
  assign n4534 = n4533 ^ n4532 ;
  assign n4535 = n4534 ^ n4515 ;
  assign n4536 = n4527 & ~n4535 ;
  assign n4537 = n4536 ^ n4533 ;
  assign n4538 = n4537 ^ n2527 ;
  assign n4540 = n4538 ^ x240 ;
  assign n4539 = n4538 ^ n4521 ;
  assign n4541 = n4540 ^ n4539 ;
  assign n4542 = ~n4526 & n4541 ;
  assign n4543 = n4542 ^ n4540 ;
  assign n4697 = n4543 ^ x255 ;
  assign n4698 = ~n4696 & n4697 ;
  assign n4553 = n4532 ^ n2527 ;
  assign n4554 = ~n4537 & n4553 ;
  assign n4555 = n4554 ^ n2527 ;
  assign n4556 = n4555 ^ n3295 ;
  assign n4544 = n3997 ^ n3996 ;
  assign n4545 = n4544 ^ n3623 ;
  assign n4546 = n4545 ^ n4186 ;
  assign n4547 = n4546 ^ n4544 ;
  assign n4548 = ~n4187 & ~n4547 ;
  assign n4549 = n4548 ^ n4545 ;
  assign n4550 = n4549 ^ n3302 ;
  assign n4551 = ~n3770 & ~n4550 ;
  assign n4552 = n4551 ^ n3302 ;
  assign n4557 = n4556 ^ n4552 ;
  assign n4559 = n4557 ^ x255 ;
  assign n4558 = n4557 ^ n4538 ;
  assign n4560 = n4559 ^ n4558 ;
  assign n4561 = n4543 & ~n4560 ;
  assign n4562 = n4561 ^ n4559 ;
  assign n4699 = n4562 ^ x254 ;
  assign n4700 = ~n4698 & ~n4699 ;
  assign n4563 = n4555 ^ n4552 ;
  assign n4564 = n3785 ^ n3352 ;
  assign n4566 = n4544 ^ n3771 ;
  assign n4567 = n4549 & n4566 ;
  assign n4568 = n4567 ^ n3771 ;
  assign n4565 = n3999 ^ n3998 ;
  assign n4569 = n4568 ^ n4565 ;
  assign n4570 = n4569 ^ n3785 ;
  assign n4571 = ~n4564 & n4570 ;
  assign n4572 = n4571 ^ n3352 ;
  assign n4573 = n4572 ^ n3295 ;
  assign n4574 = n4573 ^ n4552 ;
  assign n4575 = n4574 ^ n4572 ;
  assign n4576 = ~n4563 & n4575 ;
  assign n4577 = n4576 ^ n4573 ;
  assign n4578 = n4577 ^ n2580 ;
  assign n4580 = n4578 ^ x254 ;
  assign n4579 = n4578 ^ n4557 ;
  assign n4581 = n4580 ^ n4579 ;
  assign n4582 = n4562 & ~n4581 ;
  assign n4583 = n4582 ^ n4580 ;
  assign n4701 = n4583 ^ x253 ;
  assign n4702 = ~n4700 & n4701 ;
  assign n4588 = n3799 ^ n3391 ;
  assign n4594 = n4001 ^ n4000 ;
  assign n4590 = n3799 ^ n3785 ;
  assign n4589 = n4568 ^ n3799 ;
  assign n4591 = n4590 ^ n4589 ;
  assign n4592 = n4569 & ~n4591 ;
  assign n4593 = n4592 ^ n4590 ;
  assign n4595 = n4594 ^ n4593 ;
  assign n4596 = n4588 & ~n4595 ;
  assign n4597 = n4596 ^ n3391 ;
  assign n4584 = n4572 ^ n2580 ;
  assign n4585 = n4577 & n4584 ;
  assign n4586 = n4585 ^ n2580 ;
  assign n4587 = n4586 ^ n2618 ;
  assign n4598 = n4597 ^ n4587 ;
  assign n4600 = n4598 ^ x253 ;
  assign n4599 = n4598 ^ n4578 ;
  assign n4601 = n4600 ^ n4599 ;
  assign n4602 = n4583 & ~n4601 ;
  assign n4603 = n4602 ^ n4600 ;
  assign n4703 = n4603 ^ x252 ;
  assign n4704 = n4702 & n4703 ;
  assign n4609 = n3814 ^ n3455 ;
  assign n4615 = n4003 ^ n4002 ;
  assign n4611 = n3814 ^ n3799 ;
  assign n4610 = n4594 ^ n3814 ;
  assign n4612 = n4611 ^ n4610 ;
  assign n4613 = n4593 & n4612 ;
  assign n4614 = n4613 ^ n4611 ;
  assign n4616 = n4615 ^ n4614 ;
  assign n4617 = ~n4609 & n4616 ;
  assign n4618 = n4617 ^ n3455 ;
  assign n4604 = n4597 ^ n4586 ;
  assign n4605 = n4597 ^ n2618 ;
  assign n4606 = n4604 & ~n4605 ;
  assign n4607 = n4606 ^ n2618 ;
  assign n4608 = n4607 ^ n2665 ;
  assign n4619 = n4618 ^ n4608 ;
  assign n4621 = n4619 ^ x252 ;
  assign n4620 = n4619 ^ n4598 ;
  assign n4622 = n4621 ^ n4620 ;
  assign n4623 = n4603 & ~n4622 ;
  assign n4624 = n4623 ^ n4621 ;
  assign n4705 = n4624 ^ x251 ;
  assign n4706 = n4704 & ~n4705 ;
  assign n4630 = n3967 ^ n3483 ;
  assign n4636 = n4005 ^ n4004 ;
  assign n4632 = n3967 ^ n3814 ;
  assign n4631 = n4615 ^ n3967 ;
  assign n4633 = n4632 ^ n4631 ;
  assign n4634 = n4614 & ~n4633 ;
  assign n4635 = n4634 ^ n4632 ;
  assign n4637 = n4636 ^ n4635 ;
  assign n4638 = ~n4630 & ~n4637 ;
  assign n4639 = n4638 ^ n3483 ;
  assign n4625 = n4618 ^ n4607 ;
  assign n4626 = n4618 ^ n2665 ;
  assign n4627 = ~n4625 & n4626 ;
  assign n4628 = n4627 ^ n2665 ;
  assign n4629 = n4628 ^ n2710 ;
  assign n4640 = n4639 ^ n4629 ;
  assign n4642 = n4640 ^ x251 ;
  assign n4641 = n4640 ^ n4619 ;
  assign n4643 = n4642 ^ n4641 ;
  assign n4644 = ~n4624 & n4643 ;
  assign n4645 = n4644 ^ n4642 ;
  assign n4646 = n4645 ^ x250 ;
  assign n4707 = n4706 ^ n4646 ;
  assign n4708 = n4707 ^ n4459 ;
  assign n4709 = n4703 ^ n4702 ;
  assign n4710 = n4709 ^ n4430 ;
  assign n4711 = n4699 ^ n4698 ;
  assign n4712 = n4711 ^ n4305 ;
  assign n4782 = n4697 ^ n4696 ;
  assign n4777 = n4695 ^ n4694 ;
  assign n4713 = n4691 ^ n4690 ;
  assign n4714 = n4713 ^ n4270 ;
  assign n4716 = n4683 ^ n4682 ;
  assign n4717 = n4716 ^ n4238 ;
  assign n4718 = n4678 ^ n4677 ;
  assign n4719 = n4718 ^ n4223 ;
  assign n4720 = n4672 ^ n4647 ;
  assign n4721 = n4720 ^ n4200 ;
  assign n4725 = n4671 ^ n4648 ;
  assign n4723 = n4039 ^ n4038 ;
  assign n4724 = ~n4722 & n4723 ;
  assign n4726 = n4725 ^ n4724 ;
  assign n4727 = n4720 ^ n4193 ;
  assign n4728 = n4727 ^ n4724 ;
  assign n4729 = n4728 ^ n4720 ;
  assign n4730 = n4726 & n4729 ;
  assign n4731 = n4730 ^ n4727 ;
  assign n4732 = n4721 & n4731 ;
  assign n4733 = n4732 ^ n4200 ;
  assign n4734 = n4733 ^ n4207 ;
  assign n4735 = n4674 ^ n4673 ;
  assign n4736 = n4735 ^ n4733 ;
  assign n4737 = ~n4734 & ~n4736 ;
  assign n4738 = n4737 ^ n4207 ;
  assign n4739 = n4738 ^ n4215 ;
  assign n4740 = n4676 ^ n4675 ;
  assign n4741 = n4740 ^ n4738 ;
  assign n4742 = n4739 & n4741 ;
  assign n4743 = n4742 ^ n4215 ;
  assign n4744 = n4743 ^ n4718 ;
  assign n4745 = ~n4719 & n4744 ;
  assign n4746 = n4745 ^ n4223 ;
  assign n4747 = n4746 ^ n4230 ;
  assign n4748 = n4681 ^ n4679 ;
  assign n4749 = n4748 ^ n4746 ;
  assign n4750 = ~n4747 & ~n4749 ;
  assign n4751 = n4750 ^ n4230 ;
  assign n4752 = n4751 ^ n4716 ;
  assign n4753 = ~n4717 & n4752 ;
  assign n4754 = n4753 ^ n4238 ;
  assign n4755 = n4754 ^ n4246 ;
  assign n4756 = n4685 ^ n4684 ;
  assign n4757 = n4756 ^ n4754 ;
  assign n4758 = n4755 & ~n4757 ;
  assign n4759 = n4758 ^ n4246 ;
  assign n4760 = n4759 ^ n4254 ;
  assign n4761 = n4687 ^ n4686 ;
  assign n4762 = n4761 ^ n4759 ;
  assign n4763 = ~n4760 & n4762 ;
  assign n4764 = n4763 ^ n4254 ;
  assign n4715 = n4689 ^ n4688 ;
  assign n4765 = n4764 ^ n4715 ;
  assign n4766 = n4764 ^ n4262 ;
  assign n4767 = n4765 & ~n4766 ;
  assign n4768 = n4767 ^ n4262 ;
  assign n4769 = n4768 ^ n4713 ;
  assign n4770 = n4714 & ~n4769 ;
  assign n4771 = n4770 ^ n4270 ;
  assign n4772 = n4771 ^ n4279 ;
  assign n4773 = n4693 ^ n4692 ;
  assign n4774 = n4773 ^ n4771 ;
  assign n4775 = n4772 & n4774 ;
  assign n4776 = n4775 ^ n4279 ;
  assign n4778 = n4777 ^ n4776 ;
  assign n4779 = n4777 ^ n4287 ;
  assign n4780 = ~n4778 & n4779 ;
  assign n4781 = n4780 ^ n4287 ;
  assign n4783 = n4782 ^ n4781 ;
  assign n4784 = n4782 ^ n4296 ;
  assign n4785 = n4783 & ~n4784 ;
  assign n4786 = n4785 ^ n4296 ;
  assign n4787 = n4786 ^ n4711 ;
  assign n4788 = ~n4712 & n4787 ;
  assign n4789 = n4788 ^ n4305 ;
  assign n4790 = n4789 ^ n4310 ;
  assign n4791 = n4701 ^ n4700 ;
  assign n4792 = n4791 ^ n4789 ;
  assign n4793 = n4790 & n4792 ;
  assign n4794 = n4793 ^ n4310 ;
  assign n4795 = n4794 ^ n4709 ;
  assign n4796 = n4710 & ~n4795 ;
  assign n4797 = n4796 ^ n4430 ;
  assign n4798 = n4797 ^ n4444 ;
  assign n4799 = n4705 ^ n4704 ;
  assign n4800 = n4799 ^ n4797 ;
  assign n4801 = n4798 & n4800 ;
  assign n4802 = n4801 ^ n4444 ;
  assign n4803 = n4802 ^ n4707 ;
  assign n4804 = n4708 & n4803 ;
  assign n4805 = n4804 ^ n4459 ;
  assign n4806 = n4805 ^ n4474 ;
  assign n4829 = ~n4646 & n4706 ;
  assign n4812 = n4112 ^ n3510 ;
  assign n4818 = n4007 ^ n4006 ;
  assign n4814 = n4112 ^ n3967 ;
  assign n4813 = n4636 ^ n4112 ;
  assign n4815 = n4814 ^ n4813 ;
  assign n4816 = ~n4635 & n4815 ;
  assign n4817 = n4816 ^ n4814 ;
  assign n4819 = n4818 ^ n4817 ;
  assign n4820 = ~n4812 & n4819 ;
  assign n4821 = n4820 ^ n3510 ;
  assign n4807 = n4639 ^ n4628 ;
  assign n4808 = n4639 ^ n2710 ;
  assign n4809 = n4807 & n4808 ;
  assign n4810 = n4809 ^ n2710 ;
  assign n4811 = n4810 ^ n2756 ;
  assign n4822 = n4821 ^ n4811 ;
  assign n4824 = n4822 ^ x250 ;
  assign n4823 = n4822 ^ n4640 ;
  assign n4825 = n4824 ^ n4823 ;
  assign n4826 = ~n4645 & n4825 ;
  assign n4827 = n4826 ^ n4824 ;
  assign n4828 = n4827 ^ x249 ;
  assign n4830 = n4829 ^ n4828 ;
  assign n4831 = n4830 ^ n4805 ;
  assign n4832 = n4806 & ~n4831 ;
  assign n4833 = n4832 ^ n4474 ;
  assign n4834 = n4833 ^ n4488 ;
  assign n4853 = n4829 ^ n4822 ;
  assign n4854 = ~n4827 & n4853 ;
  assign n4851 = n4829 ^ n4827 ;
  assign n4852 = x249 & n4851 ;
  assign n4855 = n4854 ^ n4852 ;
  assign n4841 = n4140 ^ n3538 ;
  assign n4845 = n4818 ^ n4112 ;
  assign n4846 = ~n4817 & n4845 ;
  assign n4843 = n4009 ^ n4008 ;
  assign n4842 = n4818 ^ n4140 ;
  assign n4844 = n4843 ^ n4842 ;
  assign n4847 = n4846 ^ n4844 ;
  assign n4848 = n4841 & ~n4847 ;
  assign n4838 = n2805 ^ x248 ;
  assign n4839 = n4838 ^ n3538 ;
  assign n4840 = n4839 ^ n2756 ;
  assign n4849 = n4848 ^ n4840 ;
  assign n4835 = n4821 ^ n4810 ;
  assign n4836 = n4821 ^ n2756 ;
  assign n4837 = ~n4835 & ~n4836 ;
  assign n4850 = n4849 ^ n4837 ;
  assign n4856 = n4855 ^ n4850 ;
  assign n4857 = n4856 ^ n4833 ;
  assign n4858 = ~n4834 & ~n4857 ;
  assign n4859 = n4858 ^ n4488 ;
  assign n4860 = n4859 ^ n4503 ;
  assign n5880 = n4859 ^ n4650 ;
  assign n4864 = ~n4860 & ~n5880 ;
  assign n4861 = n4650 ^ n4517 ;
  assign n4865 = n4864 ^ n4861 ;
  assign n4868 = n4530 ^ n4517 ;
  assign n4866 = n4652 ^ n4650 ;
  assign n4867 = n4866 ^ n4530 ;
  assign n4869 = n4868 ^ n4867 ;
  assign n4870 = ~n4865 & n4869 ;
  assign n4871 = n4870 ^ n4868 ;
  assign n4873 = n4872 ^ n4871 ;
  assign n4874 = n4187 & n4873 ;
  assign n4875 = n4874 ^ n3623 ;
  assign n4876 = n4875 ^ n3616 ;
  assign n5051 = n4517 ^ n3610 ;
  assign n5052 = n4866 ^ n4865 ;
  assign n5053 = ~n5051 & n5052 ;
  assign n5054 = n5053 ^ n3610 ;
  assign n5042 = n4503 ^ n3747 ;
  assign n5043 = n4650 ^ n4503 ;
  assign n5044 = n5043 ^ n4859 ;
  assign n5045 = n5042 & n5044 ;
  assign n5046 = n5045 ^ n3747 ;
  assign n4877 = n4791 ^ n4790 ;
  assign n4878 = ~n4149 & n4877 ;
  assign n4879 = n4878 ^ n3704 ;
  assign n4880 = n4879 ^ n3025 ;
  assign n4989 = n4786 ^ n4305 ;
  assign n4990 = n4989 ^ n4711 ;
  assign n4991 = ~n4124 & n4990 ;
  assign n4992 = n4991 ^ n3695 ;
  assign n4981 = n4781 ^ n4296 ;
  assign n4982 = n4981 ^ n4782 ;
  assign n4983 = ~n4098 & n4982 ;
  assign n4984 = n4983 ^ n3688 ;
  assign n4973 = n4776 ^ n4287 ;
  assign n4974 = n4973 ^ n4777 ;
  assign n4975 = n4094 & ~n4974 ;
  assign n4976 = n4975 ^ n3680 ;
  assign n4966 = n4773 ^ n4772 ;
  assign n4967 = ~n4090 & n4966 ;
  assign n4968 = n4967 ^ n3671 ;
  assign n4958 = n4768 ^ n4270 ;
  assign n4959 = n4958 ^ n4713 ;
  assign n4960 = ~n4086 & ~n4959 ;
  assign n4961 = n4960 ^ n3663 ;
  assign n4951 = n4766 ^ n4715 ;
  assign n4952 = ~n4082 & n4951 ;
  assign n4953 = n4952 ^ n3654 ;
  assign n4944 = n4761 ^ n4760 ;
  assign n4945 = n4078 & ~n4944 ;
  assign n4946 = n4945 ^ n3645 ;
  assign n4937 = n4756 ^ n4755 ;
  assign n4938 = n4074 & ~n4937 ;
  assign n4939 = n4938 ^ n3637 ;
  assign n4929 = n4751 ^ n4238 ;
  assign n4930 = n4929 ^ n4716 ;
  assign n4931 = ~n4070 & n4930 ;
  assign n4932 = n4931 ^ n3406 ;
  assign n4922 = n4748 ^ n4747 ;
  assign n4923 = n4066 & ~n4922 ;
  assign n4924 = n4923 ^ n3363 ;
  assign n4914 = n4743 ^ n4223 ;
  assign n4915 = n4914 ^ n4718 ;
  assign n4916 = ~n4061 & ~n4915 ;
  assign n4917 = n4916 ^ n3323 ;
  assign n4907 = n4740 ^ n4739 ;
  assign n4908 = n4056 & ~n4907 ;
  assign n4909 = n4908 ^ n3280 ;
  assign n4900 = n4735 ^ n4734 ;
  assign n4901 = n4052 & n4900 ;
  assign n4902 = n4901 ^ n3237 ;
  assign n4893 = n4731 ^ n4200 ;
  assign n4894 = n4047 & n4893 ;
  assign n4895 = n4894 ^ n3196 ;
  assign n4885 = n4724 ^ n4193 ;
  assign n4886 = n4885 ^ n4725 ;
  assign n4887 = ~n4043 & ~n4886 ;
  assign n4888 = n4887 ^ n3157 ;
  assign n4881 = n4722 ^ n4039 ;
  assign n4882 = ~n4038 & ~n4881 ;
  assign n4883 = n4882 ^ n4039 ;
  assign n4884 = ~n3131 & ~n4883 ;
  assign n4889 = n4888 ^ n4884 ;
  assign n4890 = n4888 ^ n2600 ;
  assign n4891 = n4889 & n4890 ;
  assign n4892 = n4891 ^ n2600 ;
  assign n4896 = n4895 ^ n4892 ;
  assign n4897 = n4895 ^ n2635 ;
  assign n4898 = ~n4896 & n4897 ;
  assign n4899 = n4898 ^ n2635 ;
  assign n4903 = n4902 ^ n4899 ;
  assign n4904 = n4902 ^ n2682 ;
  assign n4905 = n4903 & ~n4904 ;
  assign n4906 = n4905 ^ n2682 ;
  assign n4910 = n4909 ^ n4906 ;
  assign n4911 = n4909 ^ n2727 ;
  assign n4912 = n4910 & n4911 ;
  assign n4913 = n4912 ^ n2727 ;
  assign n4918 = n4917 ^ n4913 ;
  assign n4919 = n4917 ^ n2772 ;
  assign n4920 = n4918 & ~n4919 ;
  assign n4921 = n4920 ^ n2772 ;
  assign n4925 = n4924 ^ n4921 ;
  assign n4926 = n4924 ^ n2814 ;
  assign n4927 = n4925 & n4926 ;
  assign n4928 = n4927 ^ n2814 ;
  assign n4933 = n4932 ^ n4928 ;
  assign n4934 = n4932 ^ n2835 ;
  assign n4935 = n4933 & ~n4934 ;
  assign n4936 = n4935 ^ n2835 ;
  assign n4940 = n4939 ^ n4936 ;
  assign n4941 = n4939 ^ n2856 ;
  assign n4942 = ~n4940 & n4941 ;
  assign n4943 = n4942 ^ n2856 ;
  assign n4947 = n4946 ^ n4943 ;
  assign n4948 = n4946 ^ n2878 ;
  assign n4949 = n4947 & n4948 ;
  assign n4950 = n4949 ^ n2878 ;
  assign n4954 = n4953 ^ n4950 ;
  assign n4955 = n4953 ^ n2900 ;
  assign n4956 = ~n4954 & ~n4955 ;
  assign n4957 = n4956 ^ n2900 ;
  assign n4962 = n4961 ^ n4957 ;
  assign n4963 = n4961 ^ n2922 ;
  assign n4964 = n4962 & n4963 ;
  assign n4965 = n4964 ^ n2922 ;
  assign n4969 = n4968 ^ n4965 ;
  assign n4970 = n4968 ^ n2948 ;
  assign n4971 = ~n4969 & n4970 ;
  assign n4972 = n4971 ^ n2948 ;
  assign n4977 = n4976 ^ n4972 ;
  assign n4978 = n4976 ^ n2965 ;
  assign n4979 = n4977 & ~n4978 ;
  assign n4980 = n4979 ^ n2965 ;
  assign n4985 = n4984 ^ n4980 ;
  assign n4986 = n4984 ^ n2986 ;
  assign n4987 = ~n4985 & ~n4986 ;
  assign n4988 = n4987 ^ n2986 ;
  assign n4993 = n4992 ^ n4988 ;
  assign n4994 = n4879 ^ n3008 ;
  assign n4995 = n4994 ^ n4879 ;
  assign n4996 = n4995 ^ n4988 ;
  assign n4997 = n4993 & ~n4996 ;
  assign n4998 = n4997 ^ n4994 ;
  assign n4999 = ~n4880 & ~n4998 ;
  assign n5000 = n4999 ^ n3025 ;
  assign n5001 = n5000 ^ n3567 ;
  assign n5002 = n4152 ^ n3416 ;
  assign n5003 = n4794 ^ n4430 ;
  assign n5004 = n5003 ^ n4709 ;
  assign n5005 = n5002 & ~n5004 ;
  assign n5006 = n5005 ^ n3627 ;
  assign n5007 = n5006 ^ n5000 ;
  assign n5008 = ~n5001 & ~n5007 ;
  assign n5009 = n5008 ^ n3567 ;
  assign n5010 = n5009 ^ n3070 ;
  assign n5011 = n4444 ^ n3716 ;
  assign n5012 = n4799 ^ n4798 ;
  assign n5013 = n5011 & n5012 ;
  assign n5014 = n5013 ^ n3716 ;
  assign n5015 = n5014 ^ n5009 ;
  assign n5016 = ~n5010 & n5015 ;
  assign n5017 = n5016 ^ n3070 ;
  assign n5018 = n5017 ^ n3091 ;
  assign n5019 = n4459 ^ n3614 ;
  assign n5020 = n4802 ^ n4459 ;
  assign n5021 = n5020 ^ n4707 ;
  assign n5022 = ~n5019 & ~n5021 ;
  assign n5023 = n5022 ^ n3614 ;
  assign n5024 = n5023 ^ n5017 ;
  assign n5025 = n5018 & ~n5024 ;
  assign n5026 = n5025 ^ n3091 ;
  assign n5027 = n5026 ^ n3111 ;
  assign n5028 = n4830 ^ n4806 ;
  assign n5029 = ~n4167 & n5028 ;
  assign n5030 = n5029 ^ n3731 ;
  assign n5031 = n5030 ^ n5026 ;
  assign n5032 = ~n5027 & ~n5031 ;
  assign n5033 = n5032 ^ n3111 ;
  assign n5034 = n5033 ^ n3145 ;
  assign n5035 = n4488 ^ n3739 ;
  assign n5036 = n4856 ^ n4834 ;
  assign n5037 = n5035 & ~n5036 ;
  assign n5038 = n5037 ^ n3739 ;
  assign n5039 = n5038 ^ n5033 ;
  assign n5040 = n5034 & n5039 ;
  assign n5041 = n5040 ^ n3145 ;
  assign n5047 = n5046 ^ n5041 ;
  assign n5048 = n5046 ^ n3181 ;
  assign n5049 = n5047 & ~n5048 ;
  assign n5050 = n5049 ^ n3181 ;
  assign n5055 = n5054 ^ n5050 ;
  assign n5056 = n4875 ^ n3217 ;
  assign n5057 = n5056 ^ n4875 ;
  assign n5058 = n5057 ^ n5050 ;
  assign n5059 = ~n5055 & ~n5058 ;
  assign n5060 = n5059 ^ n5056 ;
  assign n5061 = n4876 & ~n5060 ;
  assign n5062 = n5061 ^ n3616 ;
  assign n5247 = n5062 ^ n3302 ;
  assign n5064 = n4872 ^ n4530 ;
  assign n5065 = n4871 & ~n5064 ;
  assign n5066 = n5065 ^ n4530 ;
  assign n5063 = n4657 ^ n4655 ;
  assign n5067 = n5066 ^ n5063 ;
  assign n5068 = n5067 ^ n3771 ;
  assign n5069 = ~n4549 & n5068 ;
  assign n5070 = n5069 ^ n3771 ;
  assign n5248 = n5247 ^ n5070 ;
  assign n5086 = n5060 ^ n3616 ;
  assign n5087 = n5086 ^ x287 ;
  assign n5090 = n5038 ^ n5034 ;
  assign n5091 = n5090 ^ x274 ;
  assign n5094 = n4883 ^ n3131 ;
  assign n5095 = x263 & n5094 ;
  assign n5092 = n4884 ^ n2600 ;
  assign n5093 = n5092 ^ n4888 ;
  assign n5096 = n5095 ^ n5093 ;
  assign n5097 = n4892 ^ n2635 ;
  assign n5098 = n5097 ^ n4895 ;
  assign n5099 = n5098 ^ x262 ;
  assign n5100 = n5099 ^ n5093 ;
  assign n5101 = n5100 ^ n5098 ;
  assign n5102 = ~n5096 & n5101 ;
  assign n5103 = n5102 ^ n5099 ;
  assign n5104 = n4899 ^ n2682 ;
  assign n5105 = n5104 ^ n4902 ;
  assign n5107 = n5105 ^ x261 ;
  assign n5106 = n5105 ^ n5098 ;
  assign n5108 = n5107 ^ n5106 ;
  assign n5109 = n5103 & ~n5108 ;
  assign n5110 = n5109 ^ n5107 ;
  assign n5111 = n4906 ^ n2727 ;
  assign n5112 = n5111 ^ n4909 ;
  assign n5114 = n5112 ^ x260 ;
  assign n5113 = n5112 ^ n5105 ;
  assign n5115 = n5114 ^ n5113 ;
  assign n5116 = ~n5110 & n5115 ;
  assign n5117 = n5116 ^ n5114 ;
  assign n5118 = n4913 ^ n2772 ;
  assign n5119 = n5118 ^ n4917 ;
  assign n5121 = n5119 ^ x259 ;
  assign n5120 = n5119 ^ n5112 ;
  assign n5122 = n5121 ^ n5120 ;
  assign n5123 = n5117 & ~n5122 ;
  assign n5124 = n5123 ^ n5121 ;
  assign n5125 = n4921 ^ n2814 ;
  assign n5126 = n5125 ^ n4924 ;
  assign n5128 = n5126 ^ x258 ;
  assign n5127 = n5126 ^ n5119 ;
  assign n5129 = n5128 ^ n5127 ;
  assign n5130 = n5124 & ~n5129 ;
  assign n5131 = n5130 ^ n5128 ;
  assign n5132 = n4928 ^ n2835 ;
  assign n5133 = n5132 ^ n4932 ;
  assign n5135 = n5133 ^ x257 ;
  assign n5134 = n5133 ^ n5126 ;
  assign n5136 = n5135 ^ n5134 ;
  assign n5137 = ~n5131 & n5136 ;
  assign n5138 = n5137 ^ n5135 ;
  assign n5139 = n4936 ^ n2856 ;
  assign n5140 = n5139 ^ n4939 ;
  assign n5142 = n5140 ^ x256 ;
  assign n5141 = n5140 ^ n5133 ;
  assign n5143 = n5142 ^ n5141 ;
  assign n5144 = ~n5138 & n5143 ;
  assign n5145 = n5144 ^ n5142 ;
  assign n5146 = n4943 ^ n2878 ;
  assign n5147 = n5146 ^ n4946 ;
  assign n5149 = n5147 ^ x271 ;
  assign n5148 = n5147 ^ n5140 ;
  assign n5150 = n5149 ^ n5148 ;
  assign n5151 = n5145 & ~n5150 ;
  assign n5152 = n5151 ^ n5149 ;
  assign n5153 = n4950 ^ n2900 ;
  assign n5154 = n5153 ^ n4953 ;
  assign n5156 = n5154 ^ x270 ;
  assign n5155 = n5154 ^ n5147 ;
  assign n5157 = n5156 ^ n5155 ;
  assign n5158 = n5152 & ~n5157 ;
  assign n5159 = n5158 ^ n5156 ;
  assign n5160 = n4957 ^ n2922 ;
  assign n5161 = n5160 ^ n4961 ;
  assign n5163 = n5161 ^ x269 ;
  assign n5162 = n5161 ^ n5154 ;
  assign n5164 = n5163 ^ n5162 ;
  assign n5165 = n5159 & ~n5164 ;
  assign n5166 = n5165 ^ n5163 ;
  assign n5167 = n4965 ^ n2948 ;
  assign n5168 = n5167 ^ n4968 ;
  assign n5170 = n5168 ^ x268 ;
  assign n5169 = n5168 ^ n5161 ;
  assign n5171 = n5170 ^ n5169 ;
  assign n5172 = n5166 & ~n5171 ;
  assign n5173 = n5172 ^ n5170 ;
  assign n5174 = n4972 ^ n2965 ;
  assign n5175 = n5174 ^ n4976 ;
  assign n5177 = n5175 ^ x267 ;
  assign n5176 = n5175 ^ n5168 ;
  assign n5178 = n5177 ^ n5176 ;
  assign n5179 = ~n5173 & n5178 ;
  assign n5180 = n5179 ^ n5177 ;
  assign n5181 = n4980 ^ n2986 ;
  assign n5182 = n5181 ^ n4984 ;
  assign n5184 = n5182 ^ x266 ;
  assign n5183 = n5182 ^ n5175 ;
  assign n5185 = n5184 ^ n5183 ;
  assign n5186 = n5180 & ~n5185 ;
  assign n5187 = n5186 ^ n5184 ;
  assign n5188 = n4988 ^ n3008 ;
  assign n5189 = n5188 ^ n4992 ;
  assign n5191 = n5189 ^ x265 ;
  assign n5190 = n5189 ^ n5182 ;
  assign n5192 = n5191 ^ n5190 ;
  assign n5193 = n5187 & ~n5192 ;
  assign n5194 = n5193 ^ n5191 ;
  assign n5195 = n4998 ^ n3025 ;
  assign n5197 = n5195 ^ x264 ;
  assign n5196 = n5195 ^ n5189 ;
  assign n5198 = n5197 ^ n5196 ;
  assign n5199 = n5194 & ~n5198 ;
  assign n5200 = n5199 ^ n5197 ;
  assign n5201 = n5006 ^ n5001 ;
  assign n5203 = n5201 ^ x279 ;
  assign n5202 = n5201 ^ n5195 ;
  assign n5204 = n5203 ^ n5202 ;
  assign n5205 = n5200 & ~n5204 ;
  assign n5206 = n5205 ^ n5203 ;
  assign n5207 = n5014 ^ n5010 ;
  assign n5209 = n5207 ^ x278 ;
  assign n5208 = n5207 ^ n5201 ;
  assign n5210 = n5209 ^ n5208 ;
  assign n5211 = ~n5206 & n5210 ;
  assign n5212 = n5211 ^ n5209 ;
  assign n5213 = n5023 ^ n5018 ;
  assign n5215 = n5213 ^ x277 ;
  assign n5214 = n5213 ^ n5207 ;
  assign n5216 = n5215 ^ n5214 ;
  assign n5217 = ~n5212 & n5216 ;
  assign n5218 = n5217 ^ n5215 ;
  assign n5219 = n5030 ^ n5027 ;
  assign n5221 = n5219 ^ x276 ;
  assign n5220 = n5219 ^ n5213 ;
  assign n5222 = n5221 ^ n5220 ;
  assign n5223 = n5218 & ~n5222 ;
  assign n5224 = n5223 ^ n5221 ;
  assign n5226 = n5090 ^ x275 ;
  assign n5225 = n5219 ^ n5090 ;
  assign n5227 = n5226 ^ n5225 ;
  assign n5228 = ~n5224 & n5227 ;
  assign n5229 = n5228 ^ n5226 ;
  assign n5230 = ~n5091 & n5229 ;
  assign n5231 = n5230 ^ x274 ;
  assign n5232 = n5231 ^ x273 ;
  assign n5233 = n5041 ^ n3181 ;
  assign n5234 = n5233 ^ n5046 ;
  assign n5235 = n5234 ^ n5231 ;
  assign n5236 = n5232 & n5235 ;
  assign n5237 = n5236 ^ x273 ;
  assign n5088 = n5050 ^ n3217 ;
  assign n5089 = n5088 ^ n5054 ;
  assign n5238 = n5237 ^ n5089 ;
  assign n5240 = n5086 ^ x272 ;
  assign n5239 = n5237 ^ n5086 ;
  assign n5241 = n5240 ^ n5239 ;
  assign n5242 = n5238 & n5241 ;
  assign n5243 = n5242 ^ n5240 ;
  assign n5244 = ~n5087 & n5243 ;
  assign n5245 = n5244 ^ x287 ;
  assign n5246 = n5245 ^ x286 ;
  assign n5339 = n5248 ^ n5246 ;
  assign n5296 = n5110 ^ x260 ;
  assign n5297 = n5117 ^ x259 ;
  assign n5298 = ~n5296 & n5297 ;
  assign n5299 = n5124 ^ x258 ;
  assign n5300 = ~n5298 & ~n5299 ;
  assign n5301 = n5131 ^ x257 ;
  assign n5302 = ~n5300 & ~n5301 ;
  assign n5303 = n5138 ^ x256 ;
  assign n5304 = n5302 & ~n5303 ;
  assign n5305 = n5145 ^ x271 ;
  assign n5306 = ~n5304 & ~n5305 ;
  assign n5307 = n5152 ^ x270 ;
  assign n5308 = n5306 & ~n5307 ;
  assign n5309 = n5159 ^ x269 ;
  assign n5310 = n5308 & ~n5309 ;
  assign n5311 = n5166 ^ x268 ;
  assign n5312 = ~n5310 & n5311 ;
  assign n5313 = n5173 ^ x267 ;
  assign n5314 = n5312 & ~n5313 ;
  assign n5315 = n5180 ^ x266 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5317 = n5187 ^ x265 ;
  assign n5318 = n5316 & ~n5317 ;
  assign n5319 = n5194 ^ x264 ;
  assign n5320 = ~n5318 & n5319 ;
  assign n5321 = n5200 ^ x279 ;
  assign n5322 = ~n5320 & ~n5321 ;
  assign n5323 = n5206 ^ x278 ;
  assign n5324 = n5322 & n5323 ;
  assign n5325 = n5212 ^ x277 ;
  assign n5326 = n5324 & n5325 ;
  assign n5327 = n5218 ^ x276 ;
  assign n5328 = n5326 & ~n5327 ;
  assign n5329 = n5224 ^ x275 ;
  assign n5330 = n5328 & n5329 ;
  assign n5331 = n5229 ^ x274 ;
  assign n5332 = n5330 & ~n5331 ;
  assign n5333 = n5235 ^ x273 ;
  assign n5334 = n5332 & ~n5333 ;
  assign n5335 = n5238 ^ x272 ;
  assign n5336 = ~n5334 & n5335 ;
  assign n5337 = n5243 ^ x287 ;
  assign n5338 = n5336 & n5337 ;
  assign n5348 = n5339 ^ n5338 ;
  assign n5488 = n5348 ^ n4723 ;
  assign n5489 = ~n4722 & n5488 ;
  assign n5490 = n5489 ^ n4723 ;
  assign n5544 = n5490 ^ n4039 ;
  assign n5545 = x295 & ~n5544 ;
  assign n5798 = n5545 ^ x294 ;
  assign n5491 = ~n4039 & n5490 ;
  assign n5542 = n5491 ^ n3157 ;
  assign n5249 = n5248 ^ n5245 ;
  assign n5250 = n5246 & ~n5249 ;
  assign n5251 = n5250 ^ x286 ;
  assign n5341 = n5251 ^ x285 ;
  assign n5081 = n4659 ^ n4658 ;
  assign n5079 = n5063 ^ n4570 ;
  assign n5076 = n4549 ^ n3771 ;
  assign n5077 = n5076 ^ n5063 ;
  assign n5078 = ~n5067 & ~n5077 ;
  assign n5080 = n5079 ^ n5078 ;
  assign n5082 = n5081 ^ n5080 ;
  assign n5083 = ~n4569 & n5082 ;
  assign n5084 = n5083 ^ n3785 ;
  assign n5071 = n5070 ^ n5062 ;
  assign n5072 = n5070 ^ n3302 ;
  assign n5073 = n5071 & ~n5072 ;
  assign n5074 = n5073 ^ n3302 ;
  assign n5075 = n5074 ^ n3352 ;
  assign n5085 = n5084 ^ n5075 ;
  assign n5342 = n5341 ^ n5085 ;
  assign n5340 = ~n5338 & n5339 ;
  assign n5351 = n5342 ^ n5340 ;
  assign n5347 = n4723 ^ n4722 ;
  assign n5349 = ~n5347 & ~n5348 ;
  assign n5350 = n5349 ^ n4886 ;
  assign n5485 = n5351 ^ n5350 ;
  assign n5486 = ~n4726 & ~n5485 ;
  assign n5487 = n5486 ^ n4193 ;
  assign n5543 = n5542 ^ n5487 ;
  assign n5799 = n5798 ^ n5543 ;
  assign n5800 = n5544 ^ x295 ;
  assign n5801 = n5799 & n5800 ;
  assign n5546 = n5545 ^ n5543 ;
  assign n5492 = n5491 ^ n5487 ;
  assign n5252 = n5251 ^ n5085 ;
  assign n5258 = n4595 ^ n3799 ;
  assign n5259 = n4661 ^ n4660 ;
  assign n5260 = n5259 ^ n4570 ;
  assign n5261 = n5260 ^ n5081 ;
  assign n5262 = n5261 ^ n5259 ;
  assign n5263 = n5080 & n5262 ;
  assign n5264 = n5263 ^ n5260 ;
  assign n5265 = n5264 ^ n4595 ;
  assign n5266 = n5258 & n5265 ;
  assign n5267 = n5266 ^ n3799 ;
  assign n5253 = n5084 ^ n5074 ;
  assign n5254 = n5084 ^ n3352 ;
  assign n5255 = ~n5253 & ~n5254 ;
  assign n5256 = n5255 ^ n3352 ;
  assign n5257 = n5256 ^ n3391 ;
  assign n5268 = n5267 ^ n5257 ;
  assign n5269 = n5268 ^ x285 ;
  assign n5270 = n5269 ^ n5085 ;
  assign n5271 = n5270 ^ n5268 ;
  assign n5272 = ~n5252 & n5271 ;
  assign n5273 = n5272 ^ n5269 ;
  assign n5344 = n5273 ^ x284 ;
  assign n5343 = n5340 & n5342 ;
  assign n5356 = n5344 ^ n5343 ;
  assign n5352 = n5351 ^ n5349 ;
  assign n5353 = ~n5350 & ~n5352 ;
  assign n5354 = n5353 ^ n4886 ;
  assign n5355 = n5354 ^ n4893 ;
  assign n5481 = n5356 ^ n5355 ;
  assign n5482 = ~n4731 & n5481 ;
  assign n5483 = n5482 ^ n4200 ;
  assign n5493 = n5483 ^ n3157 ;
  assign n5494 = n5493 ^ n5487 ;
  assign n5495 = n5494 ^ n5483 ;
  assign n5496 = ~n5492 & ~n5495 ;
  assign n5497 = n5496 ^ n5493 ;
  assign n5547 = n5497 ^ n3196 ;
  assign n5548 = n5547 ^ x294 ;
  assign n5549 = n5548 ^ n5543 ;
  assign n5550 = n5549 ^ n5547 ;
  assign n5551 = n5546 & ~n5550 ;
  assign n5552 = n5551 ^ n5548 ;
  assign n5802 = n5552 ^ x293 ;
  assign n5803 = n5801 & n5802 ;
  assign n5357 = n5356 ^ n5354 ;
  assign n5358 = ~n5355 & ~n5357 ;
  assign n5359 = n5358 ^ n4893 ;
  assign n5389 = n5359 ^ n4900 ;
  assign n5345 = ~n5343 & ~n5344 ;
  assign n5279 = n4616 ^ n3814 ;
  assign n5285 = n4663 ^ n4662 ;
  assign n5281 = n4616 ^ n4595 ;
  assign n5280 = n5259 ^ n4616 ;
  assign n5282 = n5281 ^ n5280 ;
  assign n5283 = n5264 & n5282 ;
  assign n5284 = n5283 ^ n5281 ;
  assign n5286 = n5285 ^ n5284 ;
  assign n5287 = ~n5279 & n5286 ;
  assign n5288 = n5287 ^ n3814 ;
  assign n5274 = n5267 ^ n5256 ;
  assign n5275 = n5267 ^ n3391 ;
  assign n5276 = n5274 & n5275 ;
  assign n5277 = n5276 ^ n3391 ;
  assign n5278 = n5277 ^ n3455 ;
  assign n5289 = n5288 ^ n5278 ;
  assign n5291 = n5289 ^ x284 ;
  assign n5290 = n5289 ^ n5268 ;
  assign n5292 = n5291 ^ n5290 ;
  assign n5293 = ~n5273 & n5292 ;
  assign n5294 = n5293 ^ n5291 ;
  assign n5295 = n5294 ^ x283 ;
  assign n5346 = n5345 ^ n5295 ;
  assign n5501 = n5389 ^ n5346 ;
  assign n5502 = n4736 & ~n5501 ;
  assign n5503 = n5502 ^ n4207 ;
  assign n5484 = n5483 ^ n3196 ;
  assign n5498 = n5484 & ~n5497 ;
  assign n5499 = n5498 ^ n3196 ;
  assign n5500 = n5499 ^ n3237 ;
  assign n5553 = n5503 ^ n5500 ;
  assign n5555 = n5553 ^ x293 ;
  assign n5554 = n5553 ^ n5547 ;
  assign n5556 = n5555 ^ n5554 ;
  assign n5557 = n5552 & ~n5556 ;
  assign n5558 = n5557 ^ n5555 ;
  assign n5804 = n5558 ^ x292 ;
  assign n5805 = n5803 & n5804 ;
  assign n5360 = n5359 ^ n5346 ;
  assign n5390 = n5360 & n5389 ;
  assign n5391 = n5390 ^ n4900 ;
  assign n5508 = n5391 ^ n4907 ;
  assign n5370 = n4637 ^ n3967 ;
  assign n5371 = n4665 ^ n4664 ;
  assign n5373 = n5371 ^ n4616 ;
  assign n5372 = n5371 ^ n5285 ;
  assign n5374 = n5373 ^ n5372 ;
  assign n5375 = ~n5284 & ~n5374 ;
  assign n5376 = n5375 ^ n5373 ;
  assign n5377 = n5376 ^ n4637 ;
  assign n5378 = ~n5370 & ~n5377 ;
  assign n5379 = n5378 ^ n3967 ;
  assign n5365 = n5288 ^ n5277 ;
  assign n5366 = n5288 ^ n3455 ;
  assign n5367 = ~n5365 & ~n5366 ;
  assign n5368 = n5367 ^ n3455 ;
  assign n5369 = n5368 ^ n3483 ;
  assign n5380 = n5379 ^ n5369 ;
  assign n5382 = n5380 ^ x283 ;
  assign n5381 = n5380 ^ n5289 ;
  assign n5383 = n5382 ^ n5381 ;
  assign n5384 = ~n5294 & n5383 ;
  assign n5385 = n5384 ^ n5382 ;
  assign n5386 = n5385 ^ x282 ;
  assign n5364 = n5295 & ~n5345 ;
  assign n5387 = n5386 ^ n5364 ;
  assign n5509 = n5508 ^ n5387 ;
  assign n5510 = ~n4741 & ~n5509 ;
  assign n5511 = n5510 ^ n4215 ;
  assign n5504 = n5503 ^ n5499 ;
  assign n5505 = ~n5500 & n5504 ;
  assign n5506 = n5505 ^ n3237 ;
  assign n5507 = n5506 ^ n3280 ;
  assign n5559 = n5511 ^ n5507 ;
  assign n5561 = n5559 ^ x292 ;
  assign n5560 = n5559 ^ n5553 ;
  assign n5562 = n5561 ^ n5560 ;
  assign n5563 = n5558 & ~n5562 ;
  assign n5564 = n5563 ^ n5561 ;
  assign n5806 = n5564 ^ x291 ;
  assign n5807 = ~n5805 & n5806 ;
  assign n5418 = ~n5364 & n5386 ;
  assign n5401 = n4819 ^ n4112 ;
  assign n5407 = n4667 ^ n4666 ;
  assign n5403 = n4819 ^ n4637 ;
  assign n5402 = n5371 ^ n4819 ;
  assign n5404 = n5403 ^ n5402 ;
  assign n5405 = ~n5376 & ~n5404 ;
  assign n5406 = n5405 ^ n5403 ;
  assign n5408 = n5407 ^ n5406 ;
  assign n5409 = n5401 & ~n5408 ;
  assign n5410 = n5409 ^ n4112 ;
  assign n5396 = n5379 ^ n5368 ;
  assign n5397 = n5379 ^ n3483 ;
  assign n5398 = ~n5396 & ~n5397 ;
  assign n5399 = n5398 ^ n3483 ;
  assign n5400 = n5399 ^ n3510 ;
  assign n5411 = n5410 ^ n5400 ;
  assign n5413 = n5411 ^ x282 ;
  assign n5412 = n5411 ^ n5380 ;
  assign n5414 = n5413 ^ n5412 ;
  assign n5415 = n5385 & ~n5414 ;
  assign n5416 = n5415 ^ n5413 ;
  assign n5417 = n5416 ^ x281 ;
  assign n5419 = n5418 ^ n5417 ;
  assign n5388 = n5387 ^ n4907 ;
  assign n5392 = n5391 ^ n5387 ;
  assign n5393 = ~n5388 & ~n5392 ;
  assign n5394 = n5393 ^ n4907 ;
  assign n5395 = n5394 ^ n4915 ;
  assign n5516 = n5419 ^ n5395 ;
  assign n5517 = ~n4744 & n5516 ;
  assign n5518 = n5517 ^ n4223 ;
  assign n5512 = n5511 ^ n5506 ;
  assign n5513 = n5507 & ~n5512 ;
  assign n5514 = n5513 ^ n3280 ;
  assign n5515 = n5514 ^ n3323 ;
  assign n5565 = n5518 ^ n5515 ;
  assign n5567 = n5565 ^ x291 ;
  assign n5566 = n5565 ^ n5559 ;
  assign n5568 = n5567 ^ n5566 ;
  assign n5569 = ~n5564 & n5568 ;
  assign n5570 = n5569 ^ n5567 ;
  assign n5808 = n5570 ^ x290 ;
  assign n5809 = ~n5807 & n5808 ;
  assign n5420 = n5419 ^ n5394 ;
  assign n5421 = n5395 & n5420 ;
  assign n5422 = n5421 ^ n4915 ;
  assign n5523 = n5422 ^ n4922 ;
  assign n5435 = n4847 ^ n4140 ;
  assign n5439 = n5407 ^ n4819 ;
  assign n5440 = n5406 & n5439 ;
  assign n5436 = n4847 ^ n4669 ;
  assign n5437 = n5436 ^ n4668 ;
  assign n5438 = n5437 ^ n5407 ;
  assign n5441 = n5440 ^ n5438 ;
  assign n5442 = n5435 & n5441 ;
  assign n5432 = n3510 ^ x280 ;
  assign n5433 = n5432 ^ n4841 ;
  assign n5429 = n5410 ^ n5399 ;
  assign n5430 = n5410 ^ n3510 ;
  assign n5431 = n5429 & ~n5430 ;
  assign n5434 = n5433 ^ n5431 ;
  assign n5443 = n5442 ^ n5434 ;
  assign n5424 = n5418 ^ n5411 ;
  assign n5427 = ~n5416 & n5424 ;
  assign n5423 = n5416 ^ n5411 ;
  assign n5425 = n5424 ^ n5423 ;
  assign n5426 = x281 & n5425 ;
  assign n5428 = n5427 ^ n5426 ;
  assign n5444 = n5443 ^ n5428 ;
  assign n5524 = n5523 ^ n5444 ;
  assign n5525 = n4749 & n5524 ;
  assign n5526 = n5525 ^ n4230 ;
  assign n5519 = n5518 ^ n5514 ;
  assign n5520 = ~n5515 & ~n5519 ;
  assign n5521 = n5520 ^ n3323 ;
  assign n5522 = n5521 ^ n3363 ;
  assign n5571 = n5526 ^ n5522 ;
  assign n5573 = n5571 ^ x290 ;
  assign n5572 = n5571 ^ n5565 ;
  assign n5574 = n5573 ^ n5572 ;
  assign n5575 = n5570 & ~n5574 ;
  assign n5576 = n5575 ^ n5573 ;
  assign n5810 = n5576 ^ x289 ;
  assign n5811 = ~n5809 & ~n5810 ;
  assign n5527 = n5526 ^ n5521 ;
  assign n5528 = n5522 & ~n5527 ;
  assign n5529 = n5528 ^ n3363 ;
  assign n5577 = n5529 ^ n3406 ;
  assign n5451 = n5094 ^ x263 ;
  assign n5445 = n5444 ^ n5422 ;
  assign n5446 = n4930 ^ n4922 ;
  assign n5447 = n5446 ^ n4930 ;
  assign n5448 = n5447 ^ n5422 ;
  assign n5449 = n5445 & n5448 ;
  assign n5450 = n5449 ^ n5446 ;
  assign n5477 = n5451 ^ n5450 ;
  assign n5478 = ~n4752 & ~n5477 ;
  assign n5479 = n5478 ^ n4238 ;
  assign n5578 = n5577 ^ n5479 ;
  assign n5580 = n5578 ^ x289 ;
  assign n5579 = n5578 ^ n5571 ;
  assign n5581 = n5580 ^ n5579 ;
  assign n5582 = n5576 & ~n5581 ;
  assign n5583 = n5582 ^ n5580 ;
  assign n5812 = n5583 ^ x288 ;
  assign n5813 = ~n5811 & ~n5812 ;
  assign n5480 = n5479 ^ n3406 ;
  assign n5530 = n5529 ^ n5479 ;
  assign n5531 = ~n5480 & ~n5530 ;
  assign n5532 = n5531 ^ n3406 ;
  assign n5584 = n5532 ^ n3637 ;
  assign n5457 = n5095 ^ x262 ;
  assign n5458 = n5457 ^ n5093 ;
  assign n5453 = n4937 ^ n4930 ;
  assign n5452 = n5451 ^ n4937 ;
  assign n5454 = n5453 ^ n5452 ;
  assign n5455 = ~n5450 & n5454 ;
  assign n5456 = n5455 ^ n5453 ;
  assign n5473 = n5458 ^ n5456 ;
  assign n5474 = n4757 & ~n5473 ;
  assign n5475 = n5474 ^ n4246 ;
  assign n5585 = n5584 ^ n5475 ;
  assign n5587 = n5585 ^ x288 ;
  assign n5586 = n5585 ^ n5578 ;
  assign n5588 = n5587 ^ n5586 ;
  assign n5589 = ~n5583 & n5588 ;
  assign n5590 = n5589 ^ n5587 ;
  assign n5814 = n5590 ^ x303 ;
  assign n5815 = n5813 & ~n5814 ;
  assign n5476 = n5475 ^ n3637 ;
  assign n5533 = n5532 ^ n5475 ;
  assign n5534 = n5476 & n5533 ;
  assign n5535 = n5534 ^ n3637 ;
  assign n5591 = n5535 ^ n3645 ;
  assign n5461 = n4944 ^ n4937 ;
  assign n5459 = n5458 ^ n4937 ;
  assign n5460 = ~n5456 & ~n5459 ;
  assign n5462 = n5461 ^ n5460 ;
  assign n5362 = n5103 ^ x261 ;
  assign n5469 = n5462 ^ n5362 ;
  assign n5470 = ~n4762 & ~n5469 ;
  assign n5471 = n5470 ^ n4254 ;
  assign n5592 = n5591 ^ n5471 ;
  assign n5594 = n5592 ^ x303 ;
  assign n5593 = n5592 ^ n5585 ;
  assign n5595 = n5594 ^ n5593 ;
  assign n5596 = ~n5590 & n5595 ;
  assign n5597 = n5596 ^ n5594 ;
  assign n5816 = n5597 ^ x302 ;
  assign n5817 = n5815 & n5816 ;
  assign n5472 = n5471 ^ n3645 ;
  assign n5536 = n5535 ^ n5471 ;
  assign n5537 = n5472 & n5536 ;
  assign n5538 = n5537 ^ n3645 ;
  assign n5539 = n5538 ^ n3654 ;
  assign n5465 = n5296 ^ n4951 ;
  assign n5363 = n5362 ^ n4944 ;
  assign n5463 = n5363 & ~n5462 ;
  assign n5464 = n5463 ^ n5362 ;
  assign n5466 = n5465 ^ n5464 ;
  assign n5467 = ~n4765 & n5466 ;
  assign n5468 = n5467 ^ n4262 ;
  assign n5540 = n5539 ^ n5468 ;
  assign n5599 = n5540 ^ x302 ;
  assign n5598 = n5592 ^ n5540 ;
  assign n5600 = n5599 ^ n5598 ;
  assign n5601 = n5597 & ~n5600 ;
  assign n5602 = n5601 ^ n5599 ;
  assign n5818 = n5602 ^ x301 ;
  assign n5819 = n5817 & n5818 ;
  assign n5615 = n5538 ^ n5468 ;
  assign n5616 = n5539 & n5615 ;
  assign n5617 = n5616 ^ n3654 ;
  assign n5618 = n5617 ^ n3663 ;
  assign n5611 = n5297 ^ n5296 ;
  assign n5605 = n5464 ^ n5296 ;
  assign n5606 = n4959 ^ n4951 ;
  assign n5607 = n5606 ^ n4959 ;
  assign n5608 = n5607 ^ n5464 ;
  assign n5609 = ~n5605 & ~n5608 ;
  assign n5610 = n5609 ^ n5606 ;
  assign n5612 = n5611 ^ n5610 ;
  assign n5613 = n4769 & ~n5612 ;
  assign n5614 = n5613 ^ n4270 ;
  assign n5619 = n5618 ^ n5614 ;
  assign n5541 = n5540 ^ x301 ;
  assign n5603 = ~n5541 & n5602 ;
  assign n5604 = n5603 ^ x301 ;
  assign n5620 = n5619 ^ n5604 ;
  assign n5820 = n5620 ^ x300 ;
  assign n5821 = ~n5819 & ~n5820 ;
  assign n5621 = n5604 ^ x300 ;
  assign n5622 = n5620 & n5621 ;
  assign n5623 = n5622 ^ x300 ;
  assign n5822 = n5623 ^ x299 ;
  assign n5633 = n5299 ^ n5298 ;
  assign n5629 = n4966 ^ n4959 ;
  assign n5628 = n5611 ^ n4966 ;
  assign n5630 = n5629 ^ n5628 ;
  assign n5631 = ~n5610 & ~n5630 ;
  assign n5632 = n5631 ^ n5629 ;
  assign n5634 = n5633 ^ n5632 ;
  assign n5635 = ~n4774 & ~n5634 ;
  assign n5636 = n5635 ^ n4279 ;
  assign n5624 = n5617 ^ n5614 ;
  assign n5625 = n5618 & n5624 ;
  assign n5626 = n5625 ^ n3663 ;
  assign n5627 = n5626 ^ n3671 ;
  assign n5637 = n5636 ^ n5627 ;
  assign n5823 = n5822 ^ n5637 ;
  assign n5824 = ~n5821 & n5823 ;
  assign n5638 = n5637 ^ n5623 ;
  assign n5649 = n5301 ^ n5300 ;
  assign n5645 = n4974 ^ n4966 ;
  assign n5644 = n5633 ^ n4974 ;
  assign n5646 = n5645 ^ n5644 ;
  assign n5647 = ~n5632 & n5646 ;
  assign n5648 = n5647 ^ n5645 ;
  assign n5650 = n5649 ^ n5648 ;
  assign n5651 = n4778 & n5650 ;
  assign n5652 = n5651 ^ n4287 ;
  assign n5639 = n5636 ^ n5626 ;
  assign n5640 = n5636 ^ n3671 ;
  assign n5641 = n5639 & ~n5640 ;
  assign n5642 = n5641 ^ n3671 ;
  assign n5643 = n5642 ^ n3680 ;
  assign n5653 = n5652 ^ n5643 ;
  assign n5654 = n5653 ^ x299 ;
  assign n5655 = n5654 ^ n5623 ;
  assign n5656 = n5655 ^ n5653 ;
  assign n5657 = n5638 & n5656 ;
  assign n5658 = n5657 ^ n5654 ;
  assign n5825 = n5658 ^ x298 ;
  assign n5826 = n5824 & ~n5825 ;
  assign n5669 = n5303 ^ n5302 ;
  assign n5665 = n4982 ^ n4974 ;
  assign n5664 = n5649 ^ n4982 ;
  assign n5666 = n5665 ^ n5664 ;
  assign n5667 = ~n5648 & n5666 ;
  assign n5668 = n5667 ^ n5665 ;
  assign n5670 = n5669 ^ n5668 ;
  assign n5671 = ~n4783 & ~n5670 ;
  assign n5672 = n5671 ^ n4296 ;
  assign n5659 = n5652 ^ n5642 ;
  assign n5660 = n5652 ^ n3680 ;
  assign n5661 = n5659 & n5660 ;
  assign n5662 = n5661 ^ n3680 ;
  assign n5663 = n5662 ^ n3688 ;
  assign n5673 = n5672 ^ n5663 ;
  assign n5675 = n5673 ^ x298 ;
  assign n5674 = n5673 ^ n5653 ;
  assign n5676 = n5675 ^ n5674 ;
  assign n5677 = ~n5658 & n5676 ;
  assign n5678 = n5677 ^ n5675 ;
  assign n5827 = n5678 ^ x297 ;
  assign n5828 = n5826 & ~n5827 ;
  assign n5689 = n5305 ^ n5304 ;
  assign n5685 = n4990 ^ n4982 ;
  assign n5684 = n5669 ^ n4990 ;
  assign n5686 = n5685 ^ n5684 ;
  assign n5687 = ~n5668 & n5686 ;
  assign n5688 = n5687 ^ n5685 ;
  assign n5690 = n5689 ^ n5688 ;
  assign n5691 = ~n4787 & n5690 ;
  assign n5692 = n5691 ^ n4305 ;
  assign n5679 = n5672 ^ n5662 ;
  assign n5680 = n5672 ^ n3688 ;
  assign n5681 = ~n5679 & ~n5680 ;
  assign n5682 = n5681 ^ n3688 ;
  assign n5683 = n5682 ^ n3695 ;
  assign n5693 = n5692 ^ n5683 ;
  assign n5695 = n5693 ^ x297 ;
  assign n5694 = n5693 ^ n5673 ;
  assign n5696 = n5695 ^ n5694 ;
  assign n5697 = ~n5678 & n5696 ;
  assign n5698 = n5697 ^ n5695 ;
  assign n5829 = n5698 ^ x296 ;
  assign n5830 = n5828 & n5829 ;
  assign n5706 = n5689 ^ n4990 ;
  assign n5707 = n5688 & n5706 ;
  assign n5705 = n4990 ^ n4877 ;
  assign n5708 = n5707 ^ n5705 ;
  assign n5704 = n5307 ^ n5306 ;
  assign n5709 = n5708 ^ n5704 ;
  assign n5710 = ~n4792 & ~n5709 ;
  assign n5711 = n5710 ^ n4310 ;
  assign n5699 = n5692 ^ n5682 ;
  assign n5700 = n5692 ^ n3695 ;
  assign n5701 = n5699 & ~n5700 ;
  assign n5702 = n5701 ^ n3695 ;
  assign n5703 = n5702 ^ n3704 ;
  assign n5712 = n5711 ^ n5703 ;
  assign n5714 = n5712 ^ x296 ;
  assign n5713 = n5712 ^ n5693 ;
  assign n5715 = n5714 ^ n5713 ;
  assign n5716 = n5698 & ~n5715 ;
  assign n5717 = n5716 ^ n5714 ;
  assign n5831 = n5717 ^ x311 ;
  assign n5832 = ~n5830 & ~n5831 ;
  assign n5718 = n5711 ^ n5702 ;
  assign n5720 = n5704 ^ n4877 ;
  assign n5721 = n5708 & ~n5720 ;
  assign n5722 = n5721 ^ n4877 ;
  assign n5719 = n5309 ^ n5308 ;
  assign n5723 = n5722 ^ n5719 ;
  assign n5724 = n5723 ^ n5004 ;
  assign n5725 = n4795 & n5724 ;
  assign n5726 = n5725 ^ n4430 ;
  assign n5727 = n5726 ^ n3704 ;
  assign n5728 = n5727 ^ n5726 ;
  assign n5729 = n5728 ^ n5702 ;
  assign n5730 = n5718 & n5729 ;
  assign n5731 = n5730 ^ n5727 ;
  assign n5732 = n5731 ^ n3627 ;
  assign n5734 = n5732 ^ x311 ;
  assign n5733 = n5732 ^ n5712 ;
  assign n5735 = n5734 ^ n5733 ;
  assign n5736 = n5717 & ~n5735 ;
  assign n5737 = n5736 ^ n5734 ;
  assign n5833 = n5737 ^ x310 ;
  assign n5834 = n5832 & n5833 ;
  assign n5747 = n5311 ^ n5310 ;
  assign n5743 = n5012 ^ n5004 ;
  assign n5742 = n5722 ^ n5012 ;
  assign n5744 = n5743 ^ n5742 ;
  assign n5745 = n5723 & ~n5744 ;
  assign n5746 = n5745 ^ n5743 ;
  assign n5748 = n5747 ^ n5746 ;
  assign n5749 = ~n4800 & ~n5748 ;
  assign n5750 = n5749 ^ n4444 ;
  assign n5738 = n5726 ^ n3627 ;
  assign n5739 = n5731 & n5738 ;
  assign n5740 = n5739 ^ n3627 ;
  assign n5741 = n5740 ^ n3716 ;
  assign n5751 = n5750 ^ n5741 ;
  assign n5753 = n5751 ^ x310 ;
  assign n5752 = n5751 ^ n5732 ;
  assign n5754 = n5753 ^ n5752 ;
  assign n5755 = ~n5737 & n5754 ;
  assign n5756 = n5755 ^ n5753 ;
  assign n5835 = n5756 ^ x309 ;
  assign n5836 = ~n5834 & n5835 ;
  assign n5767 = n5313 ^ n5312 ;
  assign n5763 = n5021 ^ n5012 ;
  assign n5762 = n5747 ^ n5021 ;
  assign n5764 = n5763 ^ n5762 ;
  assign n5765 = ~n5746 & n5764 ;
  assign n5766 = n5765 ^ n5763 ;
  assign n5768 = n5767 ^ n5766 ;
  assign n5769 = ~n4803 & ~n5768 ;
  assign n5770 = n5769 ^ n4459 ;
  assign n5757 = n5750 ^ n5740 ;
  assign n5758 = n5750 ^ n3716 ;
  assign n5759 = ~n5757 & n5758 ;
  assign n5760 = n5759 ^ n3716 ;
  assign n5761 = n5760 ^ n3614 ;
  assign n5771 = n5770 ^ n5761 ;
  assign n5773 = n5771 ^ x309 ;
  assign n5772 = n5771 ^ n5751 ;
  assign n5774 = n5773 ^ n5772 ;
  assign n5775 = n5756 & ~n5774 ;
  assign n5776 = n5775 ^ n5773 ;
  assign n5837 = n5776 ^ x308 ;
  assign n5838 = ~n5836 & n5837 ;
  assign n5787 = n5315 ^ n5314 ;
  assign n5783 = n5028 ^ n5021 ;
  assign n5782 = n5767 ^ n5028 ;
  assign n5784 = n5783 ^ n5782 ;
  assign n5785 = ~n5766 & ~n5784 ;
  assign n5786 = n5785 ^ n5783 ;
  assign n5788 = n5787 ^ n5786 ;
  assign n5789 = n4831 & ~n5788 ;
  assign n5790 = n5789 ^ n4474 ;
  assign n5777 = n5770 ^ n5760 ;
  assign n5778 = n5770 ^ n3614 ;
  assign n5779 = n5777 & ~n5778 ;
  assign n5780 = n5779 ^ n3614 ;
  assign n5781 = n5780 ^ n3731 ;
  assign n5791 = n5790 ^ n5781 ;
  assign n5793 = n5791 ^ x308 ;
  assign n5792 = n5791 ^ n5771 ;
  assign n5794 = n5793 ^ n5792 ;
  assign n5795 = ~n5776 & n5794 ;
  assign n5796 = n5795 ^ n5793 ;
  assign n5797 = n5796 ^ x307 ;
  assign n5839 = n5838 ^ n5797 ;
  assign n5922 = n5839 ^ n5347 ;
  assign n5923 = ~n5348 & n5922 ;
  assign n5924 = n5923 ^ n5347 ;
  assign n5925 = n4723 & ~n5924 ;
  assign n5926 = n5925 ^ n4193 ;
  assign n5863 = n5797 & n5838 ;
  assign n5852 = n5317 ^ n5316 ;
  assign n5848 = n5036 ^ n5028 ;
  assign n5847 = n5787 ^ n5036 ;
  assign n5849 = n5848 ^ n5847 ;
  assign n5850 = ~n5786 & n5849 ;
  assign n5851 = n5850 ^ n5848 ;
  assign n5853 = n5852 ^ n5851 ;
  assign n5854 = n4857 & n5853 ;
  assign n5855 = n5854 ^ n4488 ;
  assign n5842 = n5790 ^ n5780 ;
  assign n5843 = n5790 ^ n3731 ;
  assign n5844 = n5842 & ~n5843 ;
  assign n5845 = n5844 ^ n3731 ;
  assign n5846 = n5845 ^ n3739 ;
  assign n5856 = n5855 ^ n5846 ;
  assign n5858 = n5856 ^ x307 ;
  assign n5857 = n5856 ^ n5791 ;
  assign n5859 = n5858 ^ n5857 ;
  assign n5860 = ~n5796 & n5859 ;
  assign n5861 = n5860 ^ n5858 ;
  assign n5862 = n5861 ^ x306 ;
  assign n5864 = n5863 ^ n5862 ;
  assign n5361 = n5348 ^ n5347 ;
  assign n5840 = n5361 & n5839 ;
  assign n5841 = n5840 ^ n5485 ;
  assign n5927 = n5864 ^ n5841 ;
  assign n5928 = n5352 & n5927 ;
  assign n5929 = n5928 ^ n4886 ;
  assign n5930 = n5929 ^ n5925 ;
  assign n5931 = n5926 & n5930 ;
  assign n5932 = n5931 ^ n4193 ;
  assign n5933 = n5932 ^ n4200 ;
  assign n5890 = ~n5862 & n5863 ;
  assign n5877 = n5044 ^ n5036 ;
  assign n5875 = n5852 ^ n5036 ;
  assign n5876 = ~n5851 & n5875 ;
  assign n5878 = n5877 ^ n5876 ;
  assign n5874 = n5319 ^ n5318 ;
  assign n5879 = n5878 ^ n5874 ;
  assign n5881 = ~n5879 & ~n5880 ;
  assign n5882 = n5881 ^ n4503 ;
  assign n5869 = n5855 ^ n5845 ;
  assign n5870 = n5855 ^ n3739 ;
  assign n5871 = ~n5869 & n5870 ;
  assign n5872 = n5871 ^ n3739 ;
  assign n5873 = n5872 ^ n3747 ;
  assign n5883 = n5882 ^ n5873 ;
  assign n5885 = n5883 ^ x306 ;
  assign n5884 = n5883 ^ n5856 ;
  assign n5886 = n5885 ^ n5884 ;
  assign n5887 = n5861 & ~n5886 ;
  assign n5888 = n5887 ^ n5885 ;
  assign n5889 = n5888 ^ x305 ;
  assign n5891 = n5890 ^ n5889 ;
  assign n5865 = n5864 ^ n5840 ;
  assign n5866 = ~n5841 & n5865 ;
  assign n5867 = n5866 ^ n5485 ;
  assign n5868 = n5867 ^ n5481 ;
  assign n5934 = n5891 ^ n5868 ;
  assign n5935 = n5357 & ~n5934 ;
  assign n5936 = n5935 ^ n4893 ;
  assign n5937 = n5936 ^ n5932 ;
  assign n5938 = ~n5933 & ~n5937 ;
  assign n5939 = n5938 ^ n4200 ;
  assign n5940 = n5939 ^ n4207 ;
  assign n5917 = n5889 & ~n5890 ;
  assign n5901 = n5052 ^ n4517 ;
  assign n5905 = n5052 ^ n5044 ;
  assign n5903 = n5874 ^ n5044 ;
  assign n5904 = ~n5878 & n5903 ;
  assign n5906 = n5905 ^ n5904 ;
  assign n5902 = n5321 ^ n5320 ;
  assign n5907 = n5906 ^ n5902 ;
  assign n5908 = ~n5901 & n5907 ;
  assign n5909 = n5908 ^ n4517 ;
  assign n5896 = n5882 ^ n5872 ;
  assign n5897 = n5882 ^ n3747 ;
  assign n5898 = ~n5896 & n5897 ;
  assign n5899 = n5898 ^ n3747 ;
  assign n5900 = n5899 ^ n3610 ;
  assign n5910 = n5909 ^ n5900 ;
  assign n5912 = n5910 ^ x305 ;
  assign n5911 = n5910 ^ n5883 ;
  assign n5913 = n5912 ^ n5911 ;
  assign n5914 = n5888 & ~n5913 ;
  assign n5915 = n5914 ^ n5912 ;
  assign n5916 = n5915 ^ x304 ;
  assign n5918 = n5917 ^ n5916 ;
  assign n5892 = n5891 ^ n5867 ;
  assign n5893 = ~n5868 & n5892 ;
  assign n5894 = n5893 ^ n5481 ;
  assign n5895 = n5894 ^ n5501 ;
  assign n5919 = n5918 ^ n5895 ;
  assign n5920 = ~n5360 & n5919 ;
  assign n5921 = n5920 ^ n4900 ;
  assign n6311 = n5939 ^ n5921 ;
  assign n6312 = ~n5940 & n6311 ;
  assign n6313 = n6312 ^ n4207 ;
  assign n6314 = n6313 ^ n4215 ;
  assign n6078 = n5918 ^ n5894 ;
  assign n5965 = n5909 ^ n5899 ;
  assign n5966 = n4873 ^ n4530 ;
  assign n5972 = n5323 ^ n5322 ;
  assign n5969 = n5902 ^ n5052 ;
  assign n5970 = n5906 & n5969 ;
  assign n5967 = n5052 ^ n4873 ;
  assign n5971 = n5970 ^ n5967 ;
  assign n5973 = n5972 ^ n5971 ;
  assign n5974 = ~n5966 & n5973 ;
  assign n5975 = n5974 ^ n4530 ;
  assign n5976 = n5975 ^ n3610 ;
  assign n5977 = n5976 ^ n5975 ;
  assign n5978 = n5977 ^ n5899 ;
  assign n5979 = ~n5965 & ~n5978 ;
  assign n5980 = n5979 ^ n5976 ;
  assign n5981 = n5980 ^ n3623 ;
  assign n5983 = n5981 ^ x304 ;
  assign n5982 = n5981 ^ n5910 ;
  assign n5984 = n5983 ^ n5982 ;
  assign n5985 = ~n5915 & n5984 ;
  assign n5986 = n5985 ^ n5983 ;
  assign n5987 = n5986 ^ x319 ;
  assign n5964 = n5916 & ~n5917 ;
  assign n6076 = n5987 ^ n5964 ;
  assign n6079 = n6076 ^ n5501 ;
  assign n6080 = n6079 ^ n6076 ;
  assign n6081 = n6080 ^ n5894 ;
  assign n6082 = n6078 & ~n6081 ;
  assign n6083 = n6082 ^ n6079 ;
  assign n6315 = n6083 ^ n5509 ;
  assign n6316 = n5392 & ~n6315 ;
  assign n6317 = n6316 ^ n4907 ;
  assign n6318 = n6317 ^ n6313 ;
  assign n6319 = n6314 & n6318 ;
  assign n6320 = n6319 ^ n4215 ;
  assign n6321 = n6320 ^ n4223 ;
  assign n5997 = n5975 ^ n3623 ;
  assign n5998 = n5980 & n5997 ;
  assign n5999 = n5998 ^ n3623 ;
  assign n6000 = n5999 ^ n3771 ;
  assign n5990 = n5972 ^ n4873 ;
  assign n5991 = n5971 & n5990 ;
  assign n5992 = n5991 ^ n4873 ;
  assign n5989 = n5325 ^ n5324 ;
  assign n5993 = n5992 ^ n5989 ;
  assign n5994 = n5993 ^ n5076 ;
  assign n5995 = ~n5067 & n5994 ;
  assign n5996 = n5995 ^ n5076 ;
  assign n6001 = n6000 ^ n5996 ;
  assign n6003 = n6001 ^ x319 ;
  assign n6002 = n6001 ^ n5981 ;
  assign n6004 = n6003 ^ n6002 ;
  assign n6005 = ~n5986 & n6004 ;
  assign n6006 = n6005 ^ n6003 ;
  assign n6007 = n6006 ^ x318 ;
  assign n5988 = ~n5964 & ~n5987 ;
  assign n6087 = n6007 ^ n5988 ;
  assign n6077 = n6076 ^ n5509 ;
  assign n6084 = n6077 & ~n6083 ;
  assign n6085 = n6084 ^ n5509 ;
  assign n6086 = n6085 ^ n5516 ;
  assign n6322 = n6087 ^ n6086 ;
  assign n6323 = ~n5420 & ~n6322 ;
  assign n6324 = n6323 ^ n4915 ;
  assign n6325 = n6324 ^ n6320 ;
  assign n6326 = n6321 & n6325 ;
  assign n6327 = n6326 ^ n4223 ;
  assign n6328 = n6327 ^ n4230 ;
  assign n6088 = n6087 ^ n6085 ;
  assign n6089 = ~n6086 & n6088 ;
  assign n6090 = n6089 ^ n5516 ;
  assign n6329 = n6090 ^ n5524 ;
  assign n6013 = n5082 ^ n4570 ;
  assign n6019 = n5327 ^ n5326 ;
  assign n6017 = n5989 ^ n5082 ;
  assign n6014 = n5076 ^ n5067 ;
  assign n6015 = n6014 ^ n5989 ;
  assign n6016 = n5993 & n6015 ;
  assign n6018 = n6017 ^ n6016 ;
  assign n6020 = n6019 ^ n6018 ;
  assign n6021 = n6013 & ~n6020 ;
  assign n6022 = n6021 ^ n4570 ;
  assign n6009 = n5999 ^ n5996 ;
  assign n6010 = ~n6000 & ~n6009 ;
  assign n6011 = n6010 ^ n3771 ;
  assign n6012 = n6011 ^ n3785 ;
  assign n6023 = n6022 ^ n6012 ;
  assign n6025 = n6023 ^ x318 ;
  assign n6024 = n6023 ^ n6001 ;
  assign n6026 = n6025 ^ n6024 ;
  assign n6027 = ~n6006 & n6026 ;
  assign n6028 = n6027 ^ n6025 ;
  assign n6029 = n6028 ^ x317 ;
  assign n6008 = n5988 & ~n6007 ;
  assign n6091 = n6029 ^ n6008 ;
  assign n6330 = n6329 ^ n6091 ;
  assign n6331 = ~n5445 & n6330 ;
  assign n6332 = n6331 ^ n4922 ;
  assign n6333 = n6332 ^ n6327 ;
  assign n6334 = ~n6328 & n6333 ;
  assign n6335 = n6334 ^ n4230 ;
  assign n6336 = n6335 ^ n4238 ;
  assign n6337 = n5477 ^ n4930 ;
  assign n6092 = n6091 ^ n6090 ;
  assign n6093 = n6091 ^ n5524 ;
  assign n6094 = ~n6092 & n6093 ;
  assign n6095 = n6094 ^ n5524 ;
  assign n6338 = n6095 ^ n5477 ;
  assign n6040 = n6022 ^ n3785 ;
  assign n6041 = n6022 ^ n6011 ;
  assign n6042 = ~n6040 & ~n6041 ;
  assign n6043 = n6042 ^ n3785 ;
  assign n6044 = n6043 ^ n3799 ;
  assign n6031 = n5329 ^ n5328 ;
  assign n6032 = n6031 ^ n5082 ;
  assign n6033 = n6032 ^ n6019 ;
  assign n6034 = n6033 ^ n6031 ;
  assign n6035 = n6018 & ~n6034 ;
  assign n6036 = n6035 ^ n6032 ;
  assign n6037 = n6036 ^ n4595 ;
  assign n6038 = ~n5264 & n6037 ;
  assign n6039 = n6038 ^ n4595 ;
  assign n6045 = n6044 ^ n6039 ;
  assign n6047 = n6045 ^ x317 ;
  assign n6046 = n6045 ^ n6023 ;
  assign n6048 = n6047 ^ n6046 ;
  assign n6049 = n6028 & ~n6048 ;
  assign n6050 = n6049 ^ n6047 ;
  assign n6051 = n6050 ^ x316 ;
  assign n6030 = ~n6008 & ~n6029 ;
  assign n6096 = n6051 ^ n6030 ;
  assign n6339 = n6338 ^ n6096 ;
  assign n6340 = ~n6337 & ~n6339 ;
  assign n6341 = n6340 ^ n4930 ;
  assign n6342 = n6341 ^ n6335 ;
  assign n6343 = n6336 & n6342 ;
  assign n6344 = n6343 ^ n4238 ;
  assign n6345 = n6344 ^ n4246 ;
  assign n6346 = n5473 ^ n4937 ;
  assign n6097 = n6096 ^ n6095 ;
  assign n6098 = n6096 ^ n5477 ;
  assign n6099 = ~n6097 & ~n6098 ;
  assign n6100 = n6099 ^ n5477 ;
  assign n6347 = n6100 ^ n5473 ;
  assign n6057 = n5286 ^ n4616 ;
  assign n6063 = n5331 ^ n5330 ;
  assign n6059 = n5286 ^ n5265 ;
  assign n6058 = n6031 ^ n5286 ;
  assign n6060 = n6059 ^ n6058 ;
  assign n6061 = ~n6036 & n6060 ;
  assign n6062 = n6061 ^ n6059 ;
  assign n6064 = n6063 ^ n6062 ;
  assign n6065 = n6057 & ~n6064 ;
  assign n6066 = n6065 ^ n4616 ;
  assign n6053 = n6043 ^ n6039 ;
  assign n6054 = n6044 & ~n6053 ;
  assign n6055 = n6054 ^ n3799 ;
  assign n6056 = n6055 ^ n3814 ;
  assign n6067 = n6066 ^ n6056 ;
  assign n6069 = n6067 ^ x316 ;
  assign n6068 = n6067 ^ n6045 ;
  assign n6070 = n6069 ^ n6068 ;
  assign n6071 = n6050 & ~n6070 ;
  assign n6072 = n6071 ^ n6069 ;
  assign n6073 = n6072 ^ x315 ;
  assign n6052 = ~n6030 & n6051 ;
  assign n6074 = n6073 ^ n6052 ;
  assign n6348 = n6347 ^ n6074 ;
  assign n6349 = n6346 & ~n6348 ;
  assign n6350 = n6349 ^ n4937 ;
  assign n6351 = n6350 ^ n6344 ;
  assign n6352 = n6345 & ~n6351 ;
  assign n6353 = n6352 ^ n4246 ;
  assign n6354 = n6353 ^ n4254 ;
  assign n6355 = n5469 ^ n4944 ;
  assign n6116 = n5333 ^ n5332 ;
  assign n6112 = n5377 ^ n5286 ;
  assign n6111 = n6063 ^ n5377 ;
  assign n6113 = n6112 ^ n6111 ;
  assign n6114 = n6062 & ~n6113 ;
  assign n6115 = n6114 ^ n6112 ;
  assign n6117 = n6116 ^ n6115 ;
  assign n6118 = n5376 & n6117 ;
  assign n6119 = n6118 ^ n4637 ;
  assign n6106 = n6066 ^ n3814 ;
  assign n6107 = n6066 ^ n6055 ;
  assign n6108 = ~n6106 & n6107 ;
  assign n6109 = n6108 ^ n3814 ;
  assign n6110 = n6109 ^ n3967 ;
  assign n6120 = n6119 ^ n6110 ;
  assign n6122 = n6120 ^ x315 ;
  assign n6121 = n6120 ^ n6067 ;
  assign n6123 = n6122 ^ n6121 ;
  assign n6124 = ~n6072 & n6123 ;
  assign n6125 = n6124 ^ n6122 ;
  assign n6126 = n6125 ^ x314 ;
  assign n6105 = ~n6052 & n6073 ;
  assign n6127 = n6126 ^ n6105 ;
  assign n6075 = n6074 ^ n5473 ;
  assign n6101 = n6100 ^ n6074 ;
  assign n6102 = n6075 & ~n6101 ;
  assign n6103 = n6102 ^ n5473 ;
  assign n6104 = n6103 ^ n5469 ;
  assign n6356 = n6127 ^ n6104 ;
  assign n6357 = n6355 & n6356 ;
  assign n6358 = n6357 ^ n4944 ;
  assign n6359 = n6358 ^ n6353 ;
  assign n6360 = ~n6354 & ~n6359 ;
  assign n6361 = n6360 ^ n4254 ;
  assign n6362 = n6361 ^ n4262 ;
  assign n6128 = n6127 ^ n6103 ;
  assign n6129 = n6104 & n6128 ;
  assign n6130 = n6129 ^ n5469 ;
  assign n6363 = n6130 ^ n5466 ;
  assign n6153 = n6105 & n6126 ;
  assign n6136 = n5408 ^ n4819 ;
  assign n6142 = n5335 ^ n5334 ;
  assign n6138 = n5408 ^ n5377 ;
  assign n6137 = n6116 ^ n5408 ;
  assign n6139 = n6138 ^ n6137 ;
  assign n6140 = ~n6115 & n6139 ;
  assign n6141 = n6140 ^ n6138 ;
  assign n6143 = n6142 ^ n6141 ;
  assign n6144 = ~n6136 & n6143 ;
  assign n6145 = n6144 ^ n4819 ;
  assign n6131 = n6119 ^ n6109 ;
  assign n6132 = n6119 ^ n3967 ;
  assign n6133 = ~n6131 & ~n6132 ;
  assign n6134 = n6133 ^ n3967 ;
  assign n6135 = n6134 ^ n4112 ;
  assign n6146 = n6145 ^ n6135 ;
  assign n6148 = n6146 ^ x314 ;
  assign n6147 = n6146 ^ n6120 ;
  assign n6149 = n6148 ^ n6147 ;
  assign n6150 = ~n6125 & n6149 ;
  assign n6151 = n6150 ^ n6148 ;
  assign n6152 = n6151 ^ x313 ;
  assign n6154 = n6153 ^ n6152 ;
  assign n6364 = n6363 ^ n6154 ;
  assign n6365 = n5605 & ~n6364 ;
  assign n6366 = n6365 ^ n4951 ;
  assign n6367 = n6366 ^ n6361 ;
  assign n6368 = ~n6362 & ~n6367 ;
  assign n6369 = n6368 ^ n4262 ;
  assign n6370 = n6369 ^ n4270 ;
  assign n6371 = n5612 ^ n4959 ;
  assign n6155 = n6154 ^ n6130 ;
  assign n6156 = n6154 ^ n5466 ;
  assign n6157 = n6155 & n6156 ;
  assign n6158 = n6157 ^ n5466 ;
  assign n6372 = n6158 ^ n5612 ;
  assign n6176 = n6153 ^ n6146 ;
  assign n6177 = ~n6151 & ~n6176 ;
  assign n6174 = n6153 ^ n6151 ;
  assign n6175 = ~x313 & n6174 ;
  assign n6178 = n6177 ^ n6175 ;
  assign n6165 = n5441 ^ n4847 ;
  assign n6169 = n6142 ^ n5408 ;
  assign n6170 = ~n6141 & ~n6169 ;
  assign n6166 = n5337 ^ n5336 ;
  assign n6167 = n6166 ^ n5441 ;
  assign n6168 = n6167 ^ n6142 ;
  assign n6171 = n6170 ^ n6168 ;
  assign n6172 = ~n6165 & ~n6171 ;
  assign n6162 = n4112 ^ x312 ;
  assign n6163 = n6162 ^ n5435 ;
  assign n6159 = n6145 ^ n6134 ;
  assign n6160 = n6145 ^ n4112 ;
  assign n6161 = ~n6159 & n6160 ;
  assign n6164 = n6163 ^ n6161 ;
  assign n6173 = n6172 ^ n6164 ;
  assign n6179 = n6178 ^ n6173 ;
  assign n6373 = n6372 ^ n6179 ;
  assign n6374 = n6371 & ~n6373 ;
  assign n6375 = n6374 ^ n4959 ;
  assign n6376 = n6375 ^ n6369 ;
  assign n6377 = n6370 & ~n6376 ;
  assign n6378 = n6377 ^ n4270 ;
  assign n6527 = n6378 ^ n4279 ;
  assign n6379 = n5634 ^ n4966 ;
  assign n6180 = n6179 ^ n6158 ;
  assign n6181 = n6179 ^ n5612 ;
  assign n6182 = ~n6180 & ~n6181 ;
  assign n6183 = n6182 ^ n5612 ;
  assign n5963 = n5800 ^ n5634 ;
  assign n6380 = n6183 ^ n5963 ;
  assign n6381 = ~n6379 & n6380 ;
  assign n6382 = n6381 ^ n4966 ;
  assign n6528 = n6527 ^ n6382 ;
  assign n6529 = n6528 ^ x331 ;
  assign n5942 = n5924 ^ n4723 ;
  assign n5943 = x327 & ~n5942 ;
  assign n5944 = n5943 ^ x326 ;
  assign n5945 = n5929 ^ n5926 ;
  assign n5946 = n5945 ^ n5943 ;
  assign n5947 = n5944 & n5946 ;
  assign n5948 = n5947 ^ x326 ;
  assign n5949 = n5948 ^ x325 ;
  assign n5950 = n5936 ^ n5933 ;
  assign n5951 = n5950 ^ n5948 ;
  assign n5952 = n5949 & n5951 ;
  assign n5953 = n5952 ^ x325 ;
  assign n5941 = n5940 ^ n5921 ;
  assign n5954 = n5953 ^ n5941 ;
  assign n6530 = n6317 ^ n6314 ;
  assign n6531 = n6530 ^ x324 ;
  assign n6532 = n6531 ^ n5953 ;
  assign n6533 = n6532 ^ n6530 ;
  assign n6534 = n5954 & n6533 ;
  assign n6535 = n6534 ^ n6531 ;
  assign n6536 = n6324 ^ n6321 ;
  assign n6538 = n6536 ^ x323 ;
  assign n6537 = n6536 ^ n6530 ;
  assign n6539 = n6538 ^ n6537 ;
  assign n6540 = n6535 & ~n6539 ;
  assign n6541 = n6540 ^ n6538 ;
  assign n6542 = n6332 ^ n6328 ;
  assign n6544 = n6542 ^ x322 ;
  assign n6543 = n6542 ^ n6536 ;
  assign n6545 = n6544 ^ n6543 ;
  assign n6546 = n6541 & ~n6545 ;
  assign n6547 = n6546 ^ n6544 ;
  assign n6548 = n6341 ^ n6336 ;
  assign n6550 = n6548 ^ x321 ;
  assign n6549 = n6548 ^ n6542 ;
  assign n6551 = n6550 ^ n6549 ;
  assign n6552 = ~n6547 & n6551 ;
  assign n6553 = n6552 ^ n6550 ;
  assign n6554 = n6350 ^ n6345 ;
  assign n6556 = n6554 ^ x320 ;
  assign n6555 = n6554 ^ n6548 ;
  assign n6557 = n6556 ^ n6555 ;
  assign n6558 = ~n6553 & n6557 ;
  assign n6559 = n6558 ^ n6556 ;
  assign n6560 = n6358 ^ n6354 ;
  assign n6562 = n6560 ^ x335 ;
  assign n6561 = n6560 ^ n6554 ;
  assign n6563 = n6562 ^ n6561 ;
  assign n6564 = n6559 & ~n6563 ;
  assign n6565 = n6564 ^ n6562 ;
  assign n6566 = n6366 ^ n6362 ;
  assign n6568 = n6566 ^ x334 ;
  assign n6567 = n6566 ^ n6560 ;
  assign n6569 = n6568 ^ n6567 ;
  assign n6570 = ~n6565 & n6569 ;
  assign n6571 = n6570 ^ n6568 ;
  assign n6572 = n6375 ^ n6370 ;
  assign n6574 = n6572 ^ x333 ;
  assign n6573 = n6572 ^ n6566 ;
  assign n6575 = n6574 ^ n6573 ;
  assign n6576 = n6571 & ~n6575 ;
  assign n6577 = n6576 ^ n6574 ;
  assign n6579 = n6528 ^ x332 ;
  assign n6578 = n6572 ^ n6528 ;
  assign n6580 = n6579 ^ n6578 ;
  assign n6581 = n6577 & ~n6580 ;
  assign n6582 = n6581 ^ n6579 ;
  assign n6583 = n6529 & ~n6582 ;
  assign n6584 = n6583 ^ x331 ;
  assign n6383 = n6382 ^ n6378 ;
  assign n6384 = n6382 ^ n4279 ;
  assign n6385 = n6383 & ~n6384 ;
  assign n6386 = n6385 ^ n4279 ;
  assign n6525 = n6386 ^ n4287 ;
  assign n6306 = n5650 ^ n4974 ;
  assign n6184 = n6183 ^ n5634 ;
  assign n6185 = ~n5963 & ~n6184 ;
  assign n6186 = n6185 ^ n5799 ;
  assign n6307 = n6186 ^ n5650 ;
  assign n6308 = ~n6306 & ~n6307 ;
  assign n6309 = n6308 ^ n4974 ;
  assign n6526 = n6525 ^ n6309 ;
  assign n6585 = n6584 ^ n6526 ;
  assign n6391 = n5670 ^ n4982 ;
  assign n6192 = n5802 ^ n5801 ;
  assign n6190 = n5670 ^ n5650 ;
  assign n6187 = n5799 ^ n5650 ;
  assign n6188 = n6187 ^ n5800 ;
  assign n6189 = n6186 & ~n6188 ;
  assign n6191 = n6190 ^ n6189 ;
  assign n6392 = n6192 ^ n6191 ;
  assign n6393 = ~n6391 & n6392 ;
  assign n6394 = n6393 ^ n4982 ;
  assign n6310 = n6309 ^ n4287 ;
  assign n6387 = n6386 ^ n6309 ;
  assign n6388 = n6310 & ~n6387 ;
  assign n6389 = n6388 ^ n4287 ;
  assign n6390 = n6389 ^ n4296 ;
  assign n6586 = n6394 ^ n6390 ;
  assign n6587 = n6586 ^ x330 ;
  assign n6588 = n6587 ^ n6584 ;
  assign n6589 = n6588 ^ n6586 ;
  assign n6590 = n6585 & n6589 ;
  assign n6591 = n6590 ^ n6587 ;
  assign n6395 = n6394 ^ n6389 ;
  assign n6396 = n6390 & n6395 ;
  assign n6397 = n6396 ^ n4296 ;
  assign n6522 = n6397 ^ n4305 ;
  assign n6398 = n5690 ^ n4990 ;
  assign n6199 = n5804 ^ n5803 ;
  assign n6195 = n5690 ^ n5670 ;
  assign n6193 = n6192 ^ n5670 ;
  assign n6194 = ~n6191 & n6193 ;
  assign n6196 = n6195 ^ n6194 ;
  assign n6399 = n6199 ^ n6196 ;
  assign n6400 = n6398 & n6399 ;
  assign n6401 = n6400 ^ n4990 ;
  assign n6523 = n6522 ^ n6401 ;
  assign n6593 = n6523 ^ x329 ;
  assign n6592 = n6586 ^ n6523 ;
  assign n6594 = n6593 ^ n6592 ;
  assign n6595 = ~n6591 & n6594 ;
  assign n6596 = n6595 ^ n6593 ;
  assign n6718 = n6596 ^ x328 ;
  assign n5955 = n5954 ^ x324 ;
  assign n5956 = n5942 ^ x327 ;
  assign n5957 = n5946 ^ x326 ;
  assign n5958 = ~n5956 & ~n5957 ;
  assign n5959 = n5951 ^ x325 ;
  assign n5960 = n5958 & ~n5959 ;
  assign n6695 = ~n5955 & n5960 ;
  assign n6696 = n6535 ^ x323 ;
  assign n6697 = ~n6695 & n6696 ;
  assign n6698 = n6541 ^ x322 ;
  assign n6699 = n6697 & n6698 ;
  assign n6700 = n6547 ^ x321 ;
  assign n6701 = ~n6699 & n6700 ;
  assign n6702 = n6553 ^ x320 ;
  assign n6703 = ~n6701 & ~n6702 ;
  assign n6704 = n6559 ^ x335 ;
  assign n6705 = n6703 & n6704 ;
  assign n6706 = n6565 ^ x334 ;
  assign n6707 = n6705 & ~n6706 ;
  assign n6708 = n6571 ^ x333 ;
  assign n6709 = ~n6707 & ~n6708 ;
  assign n6710 = n6577 ^ x332 ;
  assign n6711 = ~n6709 & n6710 ;
  assign n6712 = n6582 ^ x331 ;
  assign n6713 = n6711 & ~n6712 ;
  assign n6714 = n6585 ^ x330 ;
  assign n6715 = ~n6713 & ~n6714 ;
  assign n6716 = n6591 ^ x329 ;
  assign n6717 = ~n6715 & ~n6716 ;
  assign n6764 = n6718 ^ n6717 ;
  assign n6880 = n6764 ^ n5361 ;
  assign n6881 = n5839 & n6880 ;
  assign n6882 = n6881 ^ n5361 ;
  assign n6985 = n6882 ^ n5347 ;
  assign n6986 = x359 & ~n6985 ;
  assign n6524 = n6523 ^ x328 ;
  assign n6597 = n6524 & ~n6596 ;
  assign n6598 = n6597 ^ x328 ;
  assign n6406 = n5709 ^ n4877 ;
  assign n6204 = n5806 ^ n5805 ;
  assign n6197 = n5709 ^ n5690 ;
  assign n6198 = n6197 ^ n5709 ;
  assign n6200 = n6199 ^ n6198 ;
  assign n6201 = ~n6196 & ~n6200 ;
  assign n6202 = n6201 ^ n6197 ;
  assign n6407 = n6204 ^ n6202 ;
  assign n6408 = ~n6406 & n6407 ;
  assign n6409 = n6408 ^ n4877 ;
  assign n6520 = n6409 ^ n4310 ;
  assign n6402 = n6401 ^ n6397 ;
  assign n6403 = n6401 ^ n4305 ;
  assign n6404 = n6402 & ~n6403 ;
  assign n6405 = n6404 ^ n4305 ;
  assign n6521 = n6520 ^ n6405 ;
  assign n6599 = n6598 ^ n6521 ;
  assign n6720 = n6599 ^ x343 ;
  assign n6719 = ~n6717 & n6718 ;
  assign n6767 = n6720 ^ n6719 ;
  assign n6763 = n5839 ^ n5361 ;
  assign n6765 = n6763 & ~n6764 ;
  assign n6766 = n6765 ^ n5927 ;
  assign n6885 = n6767 ^ n6766 ;
  assign n6886 = ~n5865 & ~n6885 ;
  assign n6887 = n6886 ^ n5485 ;
  assign n6883 = ~n5347 & n6882 ;
  assign n6884 = n6883 ^ n4886 ;
  assign n6984 = n6887 ^ n6884 ;
  assign n6987 = n6986 ^ n6984 ;
  assign n6410 = n6409 ^ n6405 ;
  assign n6203 = n5808 ^ n5807 ;
  assign n6206 = n6203 ^ n5709 ;
  assign n6205 = n6204 ^ n6203 ;
  assign n6207 = n6206 ^ n6205 ;
  assign n6208 = ~n6202 & n6207 ;
  assign n6209 = n6208 ^ n6206 ;
  assign n6302 = n6209 ^ n5004 ;
  assign n6303 = ~n5723 & ~n6302 ;
  assign n6304 = n6303 ^ n5004 ;
  assign n6411 = n6304 ^ n4310 ;
  assign n6412 = n6411 ^ n6304 ;
  assign n6413 = n6412 ^ n6405 ;
  assign n6414 = n6410 & n6413 ;
  assign n6415 = n6414 ^ n6411 ;
  assign n6600 = n6415 ^ n4430 ;
  assign n6601 = n6600 ^ x343 ;
  assign n6602 = n6601 ^ n6598 ;
  assign n6603 = n6602 ^ n6600 ;
  assign n6604 = ~n6599 & n6603 ;
  assign n6605 = n6604 ^ n6601 ;
  assign n6722 = n6605 ^ x342 ;
  assign n6721 = ~n6719 & ~n6720 ;
  assign n6772 = n6722 ^ n6721 ;
  assign n6768 = n6767 ^ n6765 ;
  assign n6769 = n6766 & n6768 ;
  assign n6770 = n6769 ^ n5927 ;
  assign n6771 = n6770 ^ n5934 ;
  assign n6892 = n6772 ^ n6771 ;
  assign n6893 = ~n5892 & n6892 ;
  assign n6894 = n6893 ^ n5481 ;
  assign n6888 = n6887 ^ n6883 ;
  assign n6889 = ~n6884 & n6888 ;
  assign n6890 = n6889 ^ n4886 ;
  assign n6891 = n6890 ^ n4893 ;
  assign n6988 = n6894 ^ n6891 ;
  assign n6989 = n6988 ^ x358 ;
  assign n6990 = n6989 ^ n6984 ;
  assign n6991 = n6990 ^ n6988 ;
  assign n6992 = ~n6987 & n6991 ;
  assign n6993 = n6992 ^ n6989 ;
  assign n6773 = n6772 ^ n6770 ;
  assign n6774 = ~n6771 & n6773 ;
  assign n6775 = n6774 ^ n5934 ;
  assign n6899 = n6775 ^ n5919 ;
  assign n6305 = n6304 ^ n4430 ;
  assign n6416 = n6305 & ~n6415 ;
  assign n6417 = n6416 ^ n4430 ;
  assign n6606 = n6417 ^ n4444 ;
  assign n6418 = n5748 ^ n5012 ;
  assign n6215 = n5810 ^ n5809 ;
  assign n6211 = n5748 ^ n5724 ;
  assign n6210 = n6203 ^ n5748 ;
  assign n6212 = n6211 ^ n6210 ;
  assign n6213 = n6209 & n6212 ;
  assign n6214 = n6213 ^ n6211 ;
  assign n6419 = n6215 ^ n6214 ;
  assign n6420 = ~n6418 & ~n6419 ;
  assign n6421 = n6420 ^ n5012 ;
  assign n6607 = n6606 ^ n6421 ;
  assign n6609 = n6607 ^ x342 ;
  assign n6608 = n6607 ^ n6600 ;
  assign n6610 = n6609 ^ n6608 ;
  assign n6611 = n6605 & ~n6610 ;
  assign n6612 = n6611 ^ n6609 ;
  assign n6724 = n6612 ^ x341 ;
  assign n6723 = n6721 & n6722 ;
  assign n6761 = n6724 ^ n6723 ;
  assign n6900 = n6899 ^ n6761 ;
  assign n6901 = ~n6078 & ~n6900 ;
  assign n6902 = n6901 ^ n5501 ;
  assign n6895 = n6894 ^ n6890 ;
  assign n6896 = ~n6891 & n6895 ;
  assign n6897 = n6896 ^ n4893 ;
  assign n6898 = n6897 ^ n4900 ;
  assign n6994 = n6902 ^ n6898 ;
  assign n6996 = n6994 ^ x357 ;
  assign n6995 = n6994 ^ n6988 ;
  assign n6997 = n6996 ^ n6995 ;
  assign n6998 = n6993 & ~n6997 ;
  assign n6999 = n6998 ^ n6996 ;
  assign n6422 = n6421 ^ n6417 ;
  assign n6423 = n6421 ^ n4444 ;
  assign n6424 = n6422 & ~n6423 ;
  assign n6425 = n6424 ^ n4444 ;
  assign n6613 = n6425 ^ n4459 ;
  assign n6221 = n5812 ^ n5811 ;
  assign n6217 = n5768 ^ n5748 ;
  assign n6216 = n6215 ^ n5768 ;
  assign n6218 = n6217 ^ n6216 ;
  assign n6219 = ~n6214 & ~n6218 ;
  assign n6220 = n6219 ^ n6217 ;
  assign n6222 = n6221 ^ n6220 ;
  assign n6426 = n5768 ^ n5021 ;
  assign n6427 = ~n6222 & n6426 ;
  assign n6428 = n6427 ^ n5021 ;
  assign n6614 = n6613 ^ n6428 ;
  assign n6616 = n6614 ^ x341 ;
  assign n6615 = n6614 ^ n6607 ;
  assign n6617 = n6616 ^ n6615 ;
  assign n6618 = ~n6612 & n6617 ;
  assign n6619 = n6618 ^ n6616 ;
  assign n6726 = n6619 ^ x340 ;
  assign n6725 = n6723 & ~n6724 ;
  assign n6780 = n6726 ^ n6725 ;
  assign n6762 = n6761 ^ n5919 ;
  assign n6776 = n6775 ^ n6761 ;
  assign n6777 = n6762 & n6776 ;
  assign n6778 = n6777 ^ n5919 ;
  assign n6779 = n6778 ^ n6315 ;
  assign n6907 = n6780 ^ n6779 ;
  assign n6908 = n6083 & ~n6907 ;
  assign n6909 = n6908 ^ n5509 ;
  assign n6903 = n6902 ^ n6897 ;
  assign n6904 = n6898 & n6903 ;
  assign n6905 = n6904 ^ n4900 ;
  assign n6906 = n6905 ^ n4907 ;
  assign n7000 = n6909 ^ n6906 ;
  assign n7002 = n7000 ^ x356 ;
  assign n7001 = n7000 ^ n6994 ;
  assign n7003 = n7002 ^ n7001 ;
  assign n7004 = n6999 & ~n7003 ;
  assign n7005 = n7004 ^ n7002 ;
  assign n6781 = n6780 ^ n6778 ;
  assign n6782 = ~n6779 & ~n6781 ;
  assign n6783 = n6782 ^ n6315 ;
  assign n6914 = n6783 ^ n6322 ;
  assign n6429 = n6428 ^ n6425 ;
  assign n6430 = n6428 ^ n4459 ;
  assign n6431 = ~n6429 & ~n6430 ;
  assign n6432 = n6431 ^ n4459 ;
  assign n6620 = n6432 ^ n4474 ;
  assign n6433 = n5788 ^ n5028 ;
  assign n6240 = n5814 ^ n5813 ;
  assign n6236 = n5788 ^ n5768 ;
  assign n6235 = n6221 ^ n5788 ;
  assign n6237 = n6236 ^ n6235 ;
  assign n6238 = n6220 & n6237 ;
  assign n6239 = n6238 ^ n6236 ;
  assign n6434 = n6240 ^ n6239 ;
  assign n6435 = ~n6433 & n6434 ;
  assign n6436 = n6435 ^ n5028 ;
  assign n6621 = n6620 ^ n6436 ;
  assign n6623 = n6621 ^ x340 ;
  assign n6622 = n6621 ^ n6614 ;
  assign n6624 = n6623 ^ n6622 ;
  assign n6625 = ~n6619 & n6624 ;
  assign n6626 = n6625 ^ n6623 ;
  assign n6728 = n6626 ^ x339 ;
  assign n6727 = n6725 & ~n6726 ;
  assign n6759 = n6728 ^ n6727 ;
  assign n6915 = n6914 ^ n6759 ;
  assign n6916 = ~n6088 & n6915 ;
  assign n6917 = n6916 ^ n5516 ;
  assign n6910 = n6909 ^ n6905 ;
  assign n6911 = ~n6906 & n6910 ;
  assign n6912 = n6911 ^ n4907 ;
  assign n6913 = n6912 ^ n4915 ;
  assign n7006 = n6917 ^ n6913 ;
  assign n7008 = n7006 ^ x355 ;
  assign n7007 = n7006 ^ n7000 ;
  assign n7009 = n7008 ^ n7007 ;
  assign n7010 = ~n7005 & n7009 ;
  assign n7011 = n7010 ^ n7008 ;
  assign n6437 = n6436 ^ n6432 ;
  assign n6438 = n6436 ^ n4474 ;
  assign n6439 = ~n6437 & n6438 ;
  assign n6440 = n6439 ^ n4474 ;
  assign n6627 = n6440 ^ n4488 ;
  assign n6441 = n5853 ^ n5036 ;
  assign n6246 = n5816 ^ n5815 ;
  assign n6242 = n5853 ^ n5788 ;
  assign n6241 = n6240 ^ n5853 ;
  assign n6243 = n6242 ^ n6241 ;
  assign n6244 = n6239 & ~n6243 ;
  assign n6245 = n6244 ^ n6242 ;
  assign n6442 = n6246 ^ n6245 ;
  assign n6443 = ~n6441 & n6442 ;
  assign n6444 = n6443 ^ n5036 ;
  assign n6628 = n6627 ^ n6444 ;
  assign n6630 = n6628 ^ x339 ;
  assign n6629 = n6628 ^ n6621 ;
  assign n6631 = n6630 ^ n6629 ;
  assign n6632 = ~n6626 & n6631 ;
  assign n6633 = n6632 ^ n6630 ;
  assign n6730 = n6633 ^ x338 ;
  assign n6729 = n6727 & ~n6728 ;
  assign n6788 = n6730 ^ n6729 ;
  assign n6760 = n6759 ^ n6322 ;
  assign n6784 = n6783 ^ n6759 ;
  assign n6785 = ~n6760 & n6784 ;
  assign n6786 = n6785 ^ n6322 ;
  assign n6787 = n6786 ^ n6330 ;
  assign n6922 = n6788 ^ n6787 ;
  assign n6923 = n6092 & ~n6922 ;
  assign n6924 = n6923 ^ n5524 ;
  assign n6918 = n6917 ^ n6912 ;
  assign n6919 = n6913 & n6918 ;
  assign n6920 = n6919 ^ n4915 ;
  assign n6921 = n6920 ^ n4922 ;
  assign n7012 = n6924 ^ n6921 ;
  assign n7014 = n7012 ^ x354 ;
  assign n7013 = n7012 ^ n7006 ;
  assign n7015 = n7014 ^ n7013 ;
  assign n7016 = ~n7011 & n7015 ;
  assign n7017 = n7016 ^ n7014 ;
  assign n6789 = n6788 ^ n6786 ;
  assign n6790 = ~n6787 & n6789 ;
  assign n6791 = n6790 ^ n6330 ;
  assign n6929 = n6791 ^ n6339 ;
  assign n6445 = n6444 ^ n6440 ;
  assign n6446 = n6444 ^ n4488 ;
  assign n6447 = n6445 & n6446 ;
  assign n6448 = n6447 ^ n4488 ;
  assign n6634 = n6448 ^ n4503 ;
  assign n6449 = n5879 ^ n5044 ;
  assign n6252 = n5818 ^ n5817 ;
  assign n6248 = n5879 ^ n5853 ;
  assign n6247 = n6246 ^ n5879 ;
  assign n6249 = n6248 ^ n6247 ;
  assign n6250 = ~n6245 & ~n6249 ;
  assign n6251 = n6250 ^ n6248 ;
  assign n6450 = n6252 ^ n6251 ;
  assign n6451 = ~n6449 & n6450 ;
  assign n6452 = n6451 ^ n5044 ;
  assign n6635 = n6634 ^ n6452 ;
  assign n6637 = n6635 ^ x338 ;
  assign n6636 = n6635 ^ n6628 ;
  assign n6638 = n6637 ^ n6636 ;
  assign n6639 = ~n6633 & n6638 ;
  assign n6640 = n6639 ^ n6637 ;
  assign n6732 = n6640 ^ x337 ;
  assign n6731 = n6729 & ~n6730 ;
  assign n6757 = n6732 ^ n6731 ;
  assign n6930 = n6929 ^ n6757 ;
  assign n6931 = n6097 & ~n6930 ;
  assign n6932 = n6931 ^ n5477 ;
  assign n6925 = n6924 ^ n6920 ;
  assign n6926 = n6921 & n6925 ;
  assign n6927 = n6926 ^ n4922 ;
  assign n6928 = n6927 ^ n4930 ;
  assign n7018 = n6932 ^ n6928 ;
  assign n7020 = n7018 ^ x353 ;
  assign n7019 = n7018 ^ n7012 ;
  assign n7021 = n7020 ^ n7019 ;
  assign n7022 = ~n7017 & n7021 ;
  assign n7023 = n7022 ^ n7020 ;
  assign n6453 = n6452 ^ n6448 ;
  assign n6454 = n6452 ^ n4503 ;
  assign n6455 = n6453 & ~n6454 ;
  assign n6456 = n6455 ^ n4503 ;
  assign n6641 = n6456 ^ n4517 ;
  assign n6457 = n5907 ^ n5052 ;
  assign n6258 = n5820 ^ n5819 ;
  assign n6254 = n5907 ^ n5879 ;
  assign n6253 = n6252 ^ n5907 ;
  assign n6255 = n6254 ^ n6253 ;
  assign n6256 = ~n6251 & n6255 ;
  assign n6257 = n6256 ^ n6254 ;
  assign n6458 = n6258 ^ n6257 ;
  assign n6459 = n6457 & ~n6458 ;
  assign n6460 = n6459 ^ n5052 ;
  assign n6642 = n6641 ^ n6460 ;
  assign n6644 = n6642 ^ x337 ;
  assign n6643 = n6642 ^ n6635 ;
  assign n6645 = n6644 ^ n6643 ;
  assign n6646 = ~n6640 & n6645 ;
  assign n6647 = n6646 ^ n6644 ;
  assign n6734 = n6647 ^ x336 ;
  assign n6733 = n6731 & ~n6732 ;
  assign n6796 = n6734 ^ n6733 ;
  assign n6758 = n6757 ^ n6339 ;
  assign n6792 = n6791 ^ n6757 ;
  assign n6793 = ~n6758 & ~n6792 ;
  assign n6794 = n6793 ^ n6339 ;
  assign n6795 = n6794 ^ n6348 ;
  assign n6937 = n6796 ^ n6795 ;
  assign n6938 = n6101 & n6937 ;
  assign n6939 = n6938 ^ n5473 ;
  assign n6933 = n6932 ^ n6927 ;
  assign n6934 = ~n6928 & ~n6933 ;
  assign n6935 = n6934 ^ n4930 ;
  assign n6936 = n6935 ^ n4937 ;
  assign n7024 = n6939 ^ n6936 ;
  assign n7026 = n7024 ^ x352 ;
  assign n7025 = n7024 ^ n7018 ;
  assign n7027 = n7026 ^ n7025 ;
  assign n7028 = ~n7023 & n7027 ;
  assign n7029 = n7028 ^ n7026 ;
  assign n6797 = n6796 ^ n6794 ;
  assign n6798 = n6795 & n6797 ;
  assign n6799 = n6798 ^ n6348 ;
  assign n6944 = n6799 ^ n6356 ;
  assign n6461 = n6460 ^ n6456 ;
  assign n6462 = n5973 ^ n4873 ;
  assign n6260 = n5973 ^ n5907 ;
  assign n6259 = n6258 ^ n5973 ;
  assign n6261 = n6260 ^ n6259 ;
  assign n6262 = ~n6257 & n6261 ;
  assign n6263 = n6262 ^ n6260 ;
  assign n6233 = n5823 ^ n5821 ;
  assign n6463 = n6263 ^ n6233 ;
  assign n6464 = n6462 & n6463 ;
  assign n6465 = n6464 ^ n4873 ;
  assign n6466 = n6465 ^ n4517 ;
  assign n6467 = n6466 ^ n6465 ;
  assign n6468 = n6467 ^ n6456 ;
  assign n6469 = n6461 & n6468 ;
  assign n6470 = n6469 ^ n6466 ;
  assign n6648 = n6470 ^ n4530 ;
  assign n6650 = n6648 ^ x336 ;
  assign n6649 = n6648 ^ n6642 ;
  assign n6651 = n6650 ^ n6649 ;
  assign n6652 = ~n6647 & n6651 ;
  assign n6653 = n6652 ^ n6650 ;
  assign n6736 = n6653 ^ x351 ;
  assign n6735 = n6733 & ~n6734 ;
  assign n6755 = n6736 ^ n6735 ;
  assign n6945 = n6944 ^ n6755 ;
  assign n6946 = ~n6128 & ~n6945 ;
  assign n6947 = n6946 ^ n5469 ;
  assign n6940 = n6939 ^ n6935 ;
  assign n6941 = ~n6936 & n6940 ;
  assign n6942 = n6941 ^ n4937 ;
  assign n6943 = n6942 ^ n4944 ;
  assign n7030 = n6947 ^ n6943 ;
  assign n7032 = n7030 ^ x367 ;
  assign n7031 = n7030 ^ n7024 ;
  assign n7033 = n7032 ^ n7031 ;
  assign n7034 = ~n7029 & n7033 ;
  assign n7035 = n7034 ^ n7032 ;
  assign n6234 = n6233 ^ n5973 ;
  assign n6264 = n6234 & n6263 ;
  assign n6265 = n6264 ^ n5973 ;
  assign n6232 = n5825 ^ n5824 ;
  assign n6266 = n6265 ^ n6232 ;
  assign n6471 = n6266 ^ n6014 ;
  assign n6472 = n5993 & ~n6471 ;
  assign n6473 = n6472 ^ n6014 ;
  assign n6475 = n6473 ^ n4530 ;
  assign n6474 = n6473 ^ n6465 ;
  assign n6476 = n6475 ^ n6474 ;
  assign n6477 = n6470 & ~n6476 ;
  assign n6478 = n6477 ^ n6475 ;
  assign n6654 = n6478 ^ n5076 ;
  assign n6656 = n6654 ^ x351 ;
  assign n6655 = n6654 ^ n6648 ;
  assign n6657 = n6656 ^ n6655 ;
  assign n6658 = ~n6653 & n6657 ;
  assign n6659 = n6658 ^ n6656 ;
  assign n6738 = n6659 ^ x350 ;
  assign n6737 = n6735 & ~n6736 ;
  assign n6804 = n6738 ^ n6737 ;
  assign n6756 = n6755 ^ n6356 ;
  assign n6800 = n6799 ^ n6755 ;
  assign n6801 = n6756 & n6800 ;
  assign n6802 = n6801 ^ n6356 ;
  assign n6803 = n6802 ^ n6364 ;
  assign n6952 = n6804 ^ n6803 ;
  assign n6953 = ~n6155 & ~n6952 ;
  assign n6954 = n6953 ^ n5466 ;
  assign n6948 = n6947 ^ n6942 ;
  assign n6949 = n6943 & ~n6948 ;
  assign n6950 = n6949 ^ n4944 ;
  assign n6951 = n6950 ^ n4951 ;
  assign n7036 = n6954 ^ n6951 ;
  assign n7038 = n7036 ^ x366 ;
  assign n7037 = n7036 ^ n7030 ;
  assign n7039 = n7038 ^ n7037 ;
  assign n7040 = n7035 & ~n7039 ;
  assign n7041 = n7040 ^ n7038 ;
  assign n7349 = n7041 ^ x365 ;
  assign n7331 = n6986 ^ x358 ;
  assign n7332 = n7331 ^ n6984 ;
  assign n7333 = n6993 ^ x357 ;
  assign n7334 = ~n7332 & n7333 ;
  assign n7335 = n6999 ^ x356 ;
  assign n7336 = n7334 & n7335 ;
  assign n7337 = n7005 ^ x355 ;
  assign n7338 = n7336 & ~n7337 ;
  assign n7339 = n7011 ^ x354 ;
  assign n7340 = n7338 & ~n7339 ;
  assign n7341 = n7017 ^ x353 ;
  assign n7342 = ~n7340 & n7341 ;
  assign n7343 = n7023 ^ x352 ;
  assign n7344 = ~n7342 & ~n7343 ;
  assign n7345 = n7029 ^ x367 ;
  assign n7346 = n7344 & ~n7345 ;
  assign n7347 = n7035 ^ x366 ;
  assign n7348 = n7346 & n7347 ;
  assign n7396 = n7349 ^ n7348 ;
  assign n7395 = n6764 ^ n6763 ;
  assign n7974 = n7396 ^ n7395 ;
  assign n7598 = n7396 ^ n6763 ;
  assign n7599 = ~n6764 & n7598 ;
  assign n7600 = n7599 ^ n6763 ;
  assign n7737 = n7600 ^ n5361 ;
  assign n7738 = x391 & n7737 ;
  assign n7601 = n5361 & n7600 ;
  assign n7603 = n7601 ^ n5485 ;
  assign n6805 = n6804 ^ n6802 ;
  assign n6806 = ~n6803 & ~n6805 ;
  assign n6807 = n6806 ^ n6364 ;
  assign n6876 = n6807 ^ n6373 ;
  assign n6739 = n6737 & ~n6738 ;
  assign n6297 = n6020 ^ n5082 ;
  assign n6272 = n5827 ^ n5826 ;
  assign n6270 = n6232 ^ n6020 ;
  assign n6267 = n6014 ^ n5993 ;
  assign n6268 = n6267 ^ n6232 ;
  assign n6269 = n6266 & n6268 ;
  assign n6271 = n6270 ^ n6269 ;
  assign n6298 = n6272 ^ n6271 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6300 = n6299 ^ n5082 ;
  assign n6480 = n6300 ^ n5076 ;
  assign n6479 = n6473 ^ n6300 ;
  assign n6481 = n6480 ^ n6479 ;
  assign n6482 = n6478 & ~n6481 ;
  assign n6483 = n6482 ^ n6480 ;
  assign n6660 = n6483 ^ n4570 ;
  assign n6662 = n6660 ^ x350 ;
  assign n6661 = n6660 ^ n6654 ;
  assign n6663 = n6662 ^ n6661 ;
  assign n6664 = ~n6659 & n6663 ;
  assign n6665 = n6664 ^ n6662 ;
  assign n6694 = n6665 ^ x349 ;
  assign n6753 = n6739 ^ n6694 ;
  assign n6877 = n6876 ^ n6753 ;
  assign n6878 = n6180 & ~n6877 ;
  assign n6879 = n6878 ^ n5612 ;
  assign n7042 = n6879 ^ n4959 ;
  assign n6955 = n6954 ^ n6950 ;
  assign n6956 = ~n6951 & n6955 ;
  assign n6957 = n6956 ^ n4951 ;
  assign n7043 = n7042 ^ n6957 ;
  assign n7045 = n7043 ^ x365 ;
  assign n7044 = n7043 ^ n7036 ;
  assign n7046 = n7045 ^ n7044 ;
  assign n7047 = n7041 & ~n7046 ;
  assign n7048 = n7047 ^ n7045 ;
  assign n7351 = n7048 ^ x364 ;
  assign n7350 = n7348 & n7349 ;
  assign n7399 = n7351 ^ n7350 ;
  assign n7397 = ~n7395 & ~n7396 ;
  assign n7398 = n7397 ^ n6885 ;
  assign n7595 = n7399 ^ n7398 ;
  assign n7596 = ~n6768 & n7595 ;
  assign n7597 = n7596 ^ n5927 ;
  assign n7736 = n7603 ^ n7597 ;
  assign n7739 = n7738 ^ n7736 ;
  assign n7602 = n7601 ^ n7597 ;
  assign n7604 = ~n7602 & ~n7603 ;
  assign n7605 = n7604 ^ n5485 ;
  assign n7607 = n7605 ^ n5481 ;
  assign n6958 = n6957 ^ n6879 ;
  assign n6871 = n6183 ^ n5800 ;
  assign n6740 = n6694 & n6739 ;
  assign n6273 = n6272 ^ n6020 ;
  assign n6274 = ~n6271 & ~n6273 ;
  assign n6275 = n6274 ^ n6020 ;
  assign n6231 = n5829 ^ n5828 ;
  assign n6276 = n6275 ^ n6231 ;
  assign n6487 = n6276 ^ n5265 ;
  assign n6488 = n6036 & ~n6487 ;
  assign n6489 = n6488 ^ n5265 ;
  assign n6301 = n6300 ^ n4570 ;
  assign n6484 = n6301 & n6483 ;
  assign n6485 = n6484 ^ n4570 ;
  assign n6486 = n6485 ^ n4595 ;
  assign n6666 = n6489 ^ n6486 ;
  assign n6668 = n6666 ^ x349 ;
  assign n6667 = n6666 ^ n6660 ;
  assign n6669 = n6668 ^ n6667 ;
  assign n6670 = n6665 & ~n6669 ;
  assign n6671 = n6670 ^ n6668 ;
  assign n6693 = n6671 ^ x348 ;
  assign n6812 = n6740 ^ n6693 ;
  assign n6754 = n6753 ^ n6373 ;
  assign n6808 = n6807 ^ n6753 ;
  assign n6809 = n6754 & ~n6808 ;
  assign n6810 = n6809 ^ n6373 ;
  assign n6811 = n6810 ^ n6380 ;
  assign n6872 = n6812 ^ n6811 ;
  assign n6873 = ~n6871 & n6872 ;
  assign n6874 = n6873 ^ n5634 ;
  assign n6959 = n6874 ^ n4959 ;
  assign n6960 = n6959 ^ n6874 ;
  assign n6961 = n6960 ^ n6879 ;
  assign n6962 = n6958 & n6961 ;
  assign n6963 = n6962 ^ n6959 ;
  assign n7049 = n6963 ^ n4966 ;
  assign n7051 = n7049 ^ x364 ;
  assign n7050 = n7049 ^ n7043 ;
  assign n7052 = n7051 ^ n7050 ;
  assign n7053 = ~n7048 & n7052 ;
  assign n7054 = n7053 ^ n7051 ;
  assign n7353 = n7054 ^ x363 ;
  assign n7352 = ~n7350 & n7351 ;
  assign n7404 = n7353 ^ n7352 ;
  assign n7400 = n7399 ^ n7397 ;
  assign n7401 = ~n7398 & n7400 ;
  assign n7402 = n7401 ^ n6885 ;
  assign n7403 = n7402 ^ n6892 ;
  assign n7592 = n7404 ^ n7403 ;
  assign n7593 = ~n6773 & n7592 ;
  assign n7594 = n7593 ^ n5934 ;
  assign n7740 = n7607 ^ n7594 ;
  assign n7741 = n7740 ^ x390 ;
  assign n7742 = n7741 ^ n7736 ;
  assign n7743 = n7742 ^ n7740 ;
  assign n7744 = n7739 & ~n7743 ;
  assign n7745 = n7744 ^ n7741 ;
  assign n7606 = n7605 ^ n7594 ;
  assign n7608 = ~n7606 & ~n7607 ;
  assign n7609 = n7608 ^ n5481 ;
  assign n7611 = n7609 ^ n5501 ;
  assign n7405 = n7404 ^ n7402 ;
  assign n7406 = ~n7403 & ~n7405 ;
  assign n7407 = n7406 ^ n6892 ;
  assign n7588 = n7407 ^ n6900 ;
  assign n6875 = n6874 ^ n4966 ;
  assign n6964 = ~n6875 & ~n6963 ;
  assign n6965 = n6964 ^ n4966 ;
  assign n6981 = n6965 ^ n4974 ;
  assign n6813 = n6812 ^ n6810 ;
  assign n6814 = ~n6811 & ~n6813 ;
  assign n6815 = n6814 ^ n6380 ;
  assign n6966 = n6815 ^ n6307 ;
  assign n6490 = n6489 ^ n6485 ;
  assign n6491 = ~n6486 & ~n6490 ;
  assign n6492 = n6491 ^ n4595 ;
  assign n6672 = n6492 ^ n4616 ;
  assign n6493 = n6064 ^ n5286 ;
  assign n6282 = n5831 ^ n5830 ;
  assign n6280 = n6231 ^ n6064 ;
  assign n6277 = n6036 ^ n5265 ;
  assign n6278 = n6277 ^ n6231 ;
  assign n6279 = n6276 & ~n6278 ;
  assign n6281 = n6280 ^ n6279 ;
  assign n6494 = n6282 ^ n6281 ;
  assign n6495 = ~n6493 & n6494 ;
  assign n6496 = n6495 ^ n5286 ;
  assign n6673 = n6672 ^ n6496 ;
  assign n6675 = n6673 ^ x348 ;
  assign n6674 = n6673 ^ n6666 ;
  assign n6676 = n6675 ^ n6674 ;
  assign n6677 = n6671 & ~n6676 ;
  assign n6678 = n6677 ^ n6675 ;
  assign n6742 = n6678 ^ x347 ;
  assign n6741 = n6693 & n6740 ;
  assign n6816 = n6742 ^ n6741 ;
  assign n6967 = n6966 ^ n6816 ;
  assign n6968 = ~n6186 & n6967 ;
  assign n6969 = n6968 ^ n5650 ;
  assign n6982 = n6981 ^ n6969 ;
  assign n7056 = n6982 ^ x363 ;
  assign n7055 = n7049 ^ n6982 ;
  assign n7057 = n7056 ^ n7055 ;
  assign n7058 = ~n7054 & n7057 ;
  assign n7059 = n7058 ^ n7056 ;
  assign n7355 = n7059 ^ x362 ;
  assign n7354 = ~n7352 & ~n7353 ;
  assign n7393 = n7355 ^ n7354 ;
  assign n7589 = n7588 ^ n7393 ;
  assign n7590 = ~n6776 & ~n7589 ;
  assign n7591 = n7590 ^ n5919 ;
  assign n7746 = n7611 ^ n7591 ;
  assign n7748 = n7746 ^ x389 ;
  assign n7747 = n7746 ^ n7740 ;
  assign n7749 = n7748 ^ n7747 ;
  assign n7750 = ~n7745 & n7749 ;
  assign n7751 = n7750 ^ n7748 ;
  assign n7898 = n7751 ^ x388 ;
  assign n7899 = n7738 ^ x390 ;
  assign n7900 = n7899 ^ n7736 ;
  assign n7901 = n7745 ^ x389 ;
  assign n7902 = ~n7900 & n7901 ;
  assign n7903 = ~n7898 & n7902 ;
  assign n7610 = n7609 ^ n7591 ;
  assign n7612 = ~n7610 & ~n7611 ;
  assign n7613 = n7612 ^ n5501 ;
  assign n7615 = n7613 ^ n5509 ;
  assign n6983 = n6982 ^ x362 ;
  assign n7060 = ~n6983 & n7059 ;
  assign n7061 = n7060 ^ x362 ;
  assign n7357 = n7061 ^ x361 ;
  assign n6975 = n6392 ^ n5670 ;
  assign n6817 = n6816 ^ n6815 ;
  assign n6818 = n6816 ^ n6307 ;
  assign n6819 = n6817 & n6818 ;
  assign n6820 = n6819 ^ n6307 ;
  assign n6976 = n6820 ^ n6392 ;
  assign n6497 = n6496 ^ n6492 ;
  assign n6498 = n6496 ^ n4616 ;
  assign n6499 = n6497 & n6498 ;
  assign n6500 = n6499 ^ n4616 ;
  assign n6679 = n6500 ^ n4637 ;
  assign n6501 = n6117 ^ n5377 ;
  assign n6288 = n5833 ^ n5832 ;
  assign n6284 = n6117 ^ n6064 ;
  assign n6283 = n6282 ^ n6117 ;
  assign n6285 = n6284 ^ n6283 ;
  assign n6286 = n6281 & ~n6285 ;
  assign n6287 = n6286 ^ n6284 ;
  assign n6502 = n6288 ^ n6287 ;
  assign n6503 = ~n6501 & ~n6502 ;
  assign n6504 = n6503 ^ n5377 ;
  assign n6680 = n6679 ^ n6504 ;
  assign n6682 = n6680 ^ x347 ;
  assign n6681 = n6680 ^ n6673 ;
  assign n6683 = n6682 ^ n6681 ;
  assign n6684 = n6678 & ~n6683 ;
  assign n6685 = n6684 ^ n6682 ;
  assign n6744 = n6685 ^ x346 ;
  assign n6743 = n6741 & n6742 ;
  assign n6821 = n6744 ^ n6743 ;
  assign n6977 = n6976 ^ n6821 ;
  assign n6978 = ~n6975 & ~n6977 ;
  assign n6979 = n6978 ^ n5670 ;
  assign n6970 = n6969 ^ n6965 ;
  assign n6971 = n6969 ^ n4974 ;
  assign n6972 = ~n6970 & ~n6971 ;
  assign n6973 = n6972 ^ n4974 ;
  assign n6974 = n6973 ^ n4982 ;
  assign n6980 = n6979 ^ n6974 ;
  assign n7358 = n7357 ^ n6980 ;
  assign n7356 = ~n7354 & ~n7355 ;
  assign n7412 = n7358 ^ n7356 ;
  assign n7394 = n7393 ^ n6900 ;
  assign n7408 = n7407 ^ n7393 ;
  assign n7409 = ~n7394 & ~n7408 ;
  assign n7410 = n7409 ^ n6900 ;
  assign n7411 = n7410 ^ n6907 ;
  assign n7585 = n7412 ^ n7411 ;
  assign n7586 = n6781 & ~n7585 ;
  assign n7587 = n7586 ^ n6315 ;
  assign n7752 = n7615 ^ n7587 ;
  assign n7754 = n7752 ^ x388 ;
  assign n7753 = n7752 ^ n7746 ;
  assign n7755 = n7754 ^ n7753 ;
  assign n7756 = n7751 & ~n7755 ;
  assign n7757 = n7756 ^ n7754 ;
  assign n7904 = n7757 ^ x387 ;
  assign n7905 = n7903 & ~n7904 ;
  assign n7614 = n7613 ^ n7587 ;
  assign n7616 = ~n7614 & n7615 ;
  assign n7617 = n7616 ^ n5509 ;
  assign n7619 = n7617 ^ n5516 ;
  assign n7413 = n7412 ^ n7410 ;
  assign n7414 = n7411 & ~n7413 ;
  assign n7415 = n7414 ^ n6907 ;
  assign n7581 = n7415 ^ n6915 ;
  assign n7359 = ~n7356 & ~n7358 ;
  assign n7062 = n7061 ^ n6980 ;
  assign n7068 = n6399 ^ n5690 ;
  assign n6822 = n6821 ^ n6820 ;
  assign n6823 = n6821 ^ n6392 ;
  assign n6824 = n6822 & n6823 ;
  assign n6825 = n6824 ^ n6392 ;
  assign n7069 = n6825 ^ n6399 ;
  assign n6505 = n6504 ^ n6500 ;
  assign n6506 = n6504 ^ n4637 ;
  assign n6507 = n6505 & n6506 ;
  assign n6508 = n6507 ^ n4637 ;
  assign n6686 = n6508 ^ n4819 ;
  assign n6509 = n6143 ^ n5408 ;
  assign n6290 = n6143 ^ n6117 ;
  assign n6289 = n6288 ^ n6143 ;
  assign n6291 = n6290 ^ n6289 ;
  assign n6292 = ~n6287 & n6291 ;
  assign n6293 = n6292 ^ n6290 ;
  assign n6228 = n5835 ^ n5834 ;
  assign n6510 = n6293 ^ n6228 ;
  assign n6511 = ~n6509 & n6510 ;
  assign n6512 = n6511 ^ n5408 ;
  assign n6687 = n6686 ^ n6512 ;
  assign n6689 = n6687 ^ x346 ;
  assign n6688 = n6687 ^ n6680 ;
  assign n6690 = n6689 ^ n6688 ;
  assign n6691 = ~n6685 & n6690 ;
  assign n6692 = n6691 ^ n6689 ;
  assign n6826 = n6692 ^ x345 ;
  assign n6745 = n6743 & ~n6744 ;
  assign n6827 = n6826 ^ n6745 ;
  assign n7070 = n7069 ^ n6827 ;
  assign n7071 = n7068 & n7070 ;
  assign n7072 = n7071 ^ n5690 ;
  assign n7063 = n6979 ^ n6973 ;
  assign n7064 = n6979 ^ n4982 ;
  assign n7065 = ~n7063 & ~n7064 ;
  assign n7066 = n7065 ^ n4982 ;
  assign n7067 = n7066 ^ n4990 ;
  assign n7073 = n7072 ^ n7067 ;
  assign n7074 = n7073 ^ x361 ;
  assign n7075 = n7074 ^ n6980 ;
  assign n7076 = n7075 ^ n7073 ;
  assign n7077 = ~n7062 & n7076 ;
  assign n7078 = n7077 ^ n7074 ;
  assign n7330 = n7078 ^ x360 ;
  assign n7391 = n7359 ^ n7330 ;
  assign n7582 = n7581 ^ n7391 ;
  assign n7583 = ~n6784 & ~n7582 ;
  assign n7584 = n7583 ^ n6322 ;
  assign n7758 = n7619 ^ n7584 ;
  assign n7760 = n7758 ^ x387 ;
  assign n7759 = n7758 ^ n7752 ;
  assign n7761 = n7760 ^ n7759 ;
  assign n7762 = n7757 & ~n7761 ;
  assign n7763 = n7762 ^ n7760 ;
  assign n7906 = n7763 ^ x386 ;
  assign n7907 = ~n7905 & ~n7906 ;
  assign n7618 = n7617 ^ n7584 ;
  assign n7620 = ~n7618 & ~n7619 ;
  assign n7621 = n7620 ^ n5516 ;
  assign n7623 = n7621 ^ n5524 ;
  assign n7360 = ~n7330 & n7359 ;
  assign n7079 = n7072 ^ n7066 ;
  assign n7080 = n6407 ^ n5709 ;
  assign n6828 = n6827 ^ n6825 ;
  assign n6748 = n6745 ^ n6687 ;
  assign n6749 = ~n6692 & n6748 ;
  assign n6746 = n6745 ^ n6692 ;
  assign n6747 = x345 & n6746 ;
  assign n6750 = n6749 ^ n6747 ;
  assign n6516 = n4819 ^ x344 ;
  assign n6517 = n6516 ^ n6165 ;
  assign n6513 = n6512 ^ n6508 ;
  assign n6514 = n6512 ^ n4819 ;
  assign n6515 = ~n6513 & ~n6514 ;
  assign n6518 = n6517 ^ n6515 ;
  assign n6225 = n6171 ^ n5441 ;
  assign n6230 = n6228 ^ n6143 ;
  assign n6294 = n6230 & ~n6293 ;
  assign n6226 = n6171 ^ n5836 ;
  assign n6227 = n6226 ^ n5837 ;
  assign n6229 = n6228 ^ n6227 ;
  assign n6295 = n6294 ^ n6229 ;
  assign n6296 = ~n6225 & n6295 ;
  assign n6519 = n6518 ^ n6296 ;
  assign n6751 = n6750 ^ n6519 ;
  assign n6829 = n6751 ^ n6399 ;
  assign n6830 = n6829 ^ n6825 ;
  assign n6831 = n6830 ^ n6751 ;
  assign n6832 = ~n6828 & n6831 ;
  assign n6833 = n6832 ^ n6829 ;
  assign n7081 = n6833 ^ n6407 ;
  assign n7082 = ~n7080 & ~n7081 ;
  assign n7083 = n7082 ^ n5709 ;
  assign n7084 = n7083 ^ n4990 ;
  assign n7085 = n7084 ^ n7083 ;
  assign n7086 = n7085 ^ n7066 ;
  assign n7087 = ~n7079 & n7086 ;
  assign n7088 = n7087 ^ n7084 ;
  assign n7089 = n7088 ^ n4877 ;
  assign n7091 = n7089 ^ x360 ;
  assign n7090 = n7089 ^ n7073 ;
  assign n7092 = n7091 ^ n7090 ;
  assign n7093 = ~n7078 & n7092 ;
  assign n7094 = n7093 ^ n7091 ;
  assign n7329 = n7094 ^ x375 ;
  assign n7420 = n7360 ^ n7329 ;
  assign n7392 = n7391 ^ n6915 ;
  assign n7416 = n7415 ^ n7391 ;
  assign n7417 = n7392 & n7416 ;
  assign n7418 = n7417 ^ n6915 ;
  assign n7419 = n7418 ^ n6922 ;
  assign n7578 = n7420 ^ n7419 ;
  assign n7579 = ~n6789 & ~n7578 ;
  assign n7580 = n7579 ^ n6330 ;
  assign n7764 = n7623 ^ n7580 ;
  assign n7766 = n7764 ^ x386 ;
  assign n7765 = n7764 ^ n7758 ;
  assign n7767 = n7766 ^ n7765 ;
  assign n7768 = ~n7763 & n7767 ;
  assign n7769 = n7768 ^ n7766 ;
  assign n7908 = n7769 ^ x385 ;
  assign n7909 = ~n7907 & n7908 ;
  assign n7622 = n7621 ^ n7580 ;
  assign n7624 = ~n7622 & n7623 ;
  assign n7625 = n7624 ^ n5524 ;
  assign n7627 = n7625 ^ n5477 ;
  assign n7421 = n7420 ^ n7418 ;
  assign n7422 = ~n7419 & ~n7421 ;
  assign n7423 = n7422 ^ n6922 ;
  assign n7425 = n7423 ^ n6930 ;
  assign n7361 = ~n7329 & ~n7360 ;
  assign n6752 = n6751 ^ n6407 ;
  assign n6834 = ~n6752 & n6833 ;
  assign n6835 = n6834 ^ n6407 ;
  assign n7095 = n6835 ^ n5956 ;
  assign n7096 = n7095 ^ n5724 ;
  assign n7097 = ~n6209 & ~n7096 ;
  assign n7098 = n7097 ^ n5724 ;
  assign n7100 = n7098 ^ n4877 ;
  assign n7099 = n7098 ^ n7083 ;
  assign n7101 = n7100 ^ n7099 ;
  assign n7102 = n7088 & ~n7101 ;
  assign n7103 = n7102 ^ n7100 ;
  assign n7104 = n7103 ^ n5004 ;
  assign n7106 = n7104 ^ x375 ;
  assign n7105 = n7104 ^ n7089 ;
  assign n7107 = n7106 ^ n7105 ;
  assign n7108 = n7094 & ~n7107 ;
  assign n7109 = n7108 ^ n7106 ;
  assign n7328 = n7109 ^ x374 ;
  assign n7390 = n7361 ^ n7328 ;
  assign n7575 = n7425 ^ n7390 ;
  assign n7576 = n6792 & ~n7575 ;
  assign n7577 = n7576 ^ n6339 ;
  assign n7770 = n7627 ^ n7577 ;
  assign n7772 = n7770 ^ x385 ;
  assign n7771 = n7770 ^ n7764 ;
  assign n7773 = n7772 ^ n7771 ;
  assign n7774 = ~n7769 & n7773 ;
  assign n7775 = n7774 ^ n7772 ;
  assign n7910 = n7775 ^ x384 ;
  assign n7911 = n7909 & n7910 ;
  assign n7626 = n7625 ^ n7577 ;
  assign n7628 = n7626 & ~n7627 ;
  assign n7629 = n7628 ^ n5477 ;
  assign n7631 = n7629 ^ n5473 ;
  assign n7424 = n7423 ^ n7390 ;
  assign n7426 = ~n7424 & n7425 ;
  assign n7427 = n7426 ^ n6930 ;
  assign n7571 = n7427 ^ n6937 ;
  assign n7114 = n6419 ^ n5748 ;
  assign n6224 = n6209 ^ n5724 ;
  assign n6836 = n6835 ^ n6224 ;
  assign n6837 = n5957 ^ n5956 ;
  assign n6839 = n6837 ^ n5957 ;
  assign n6840 = n6839 ^ n6224 ;
  assign n6841 = n6836 & ~n6840 ;
  assign n6842 = n6841 ^ n5957 ;
  assign n7115 = n6842 ^ n6419 ;
  assign n7116 = n7114 & ~n7115 ;
  assign n7117 = n7116 ^ n5748 ;
  assign n7110 = n7098 ^ n5004 ;
  assign n7111 = ~n7103 & ~n7110 ;
  assign n7112 = n7111 ^ n5004 ;
  assign n7113 = n7112 ^ n5012 ;
  assign n7118 = n7117 ^ n7113 ;
  assign n7120 = n7118 ^ x374 ;
  assign n7119 = n7118 ^ n7104 ;
  assign n7121 = n7120 ^ n7119 ;
  assign n7122 = n7109 & ~n7121 ;
  assign n7123 = n7122 ^ n7120 ;
  assign n7363 = n7123 ^ x373 ;
  assign n7362 = ~n7328 & n7361 ;
  assign n7428 = n7363 ^ n7362 ;
  assign n7572 = n7571 ^ n7428 ;
  assign n7573 = ~n6797 & n7572 ;
  assign n7574 = n7573 ^ n6348 ;
  assign n7776 = n7631 ^ n7574 ;
  assign n7778 = n7776 ^ x384 ;
  assign n7777 = n7776 ^ n7770 ;
  assign n7779 = n7778 ^ n7777 ;
  assign n7780 = ~n7775 & n7779 ;
  assign n7781 = n7780 ^ n7778 ;
  assign n7912 = n7781 ^ x399 ;
  assign n7913 = ~n7911 & n7912 ;
  assign n7630 = n7629 ^ n7574 ;
  assign n7632 = ~n7630 & n7631 ;
  assign n7633 = n7632 ^ n5473 ;
  assign n7635 = n7633 ^ n5469 ;
  assign n7429 = n7428 ^ n7427 ;
  assign n7430 = n7428 ^ n6937 ;
  assign n7431 = ~n7429 & ~n7430 ;
  assign n7432 = n7431 ^ n6937 ;
  assign n7567 = n7432 ^ n6945 ;
  assign n7364 = ~n7362 & ~n7363 ;
  assign n7129 = n6222 ^ n5768 ;
  assign n6844 = n6419 ^ n6222 ;
  assign n6843 = n6837 ^ n6222 ;
  assign n6845 = n6844 ^ n6843 ;
  assign n6846 = ~n6842 & ~n6845 ;
  assign n6847 = n6846 ^ n6844 ;
  assign n5962 = n5959 ^ n5958 ;
  assign n7130 = n6847 ^ n5962 ;
  assign n7131 = n7129 & ~n7130 ;
  assign n7132 = n7131 ^ n5768 ;
  assign n7124 = n7117 ^ n7112 ;
  assign n7125 = n7117 ^ n5012 ;
  assign n7126 = ~n7124 & ~n7125 ;
  assign n7127 = n7126 ^ n5012 ;
  assign n7128 = n7127 ^ n5021 ;
  assign n7133 = n7132 ^ n7128 ;
  assign n7135 = n7133 ^ x373 ;
  assign n7134 = n7133 ^ n7118 ;
  assign n7136 = n7135 ^ n7134 ;
  assign n7137 = ~n7123 & n7136 ;
  assign n7138 = n7137 ^ n7135 ;
  assign n7327 = n7138 ^ x372 ;
  assign n7388 = n7364 ^ n7327 ;
  assign n7568 = n7567 ^ n7388 ;
  assign n7569 = ~n6800 & ~n7568 ;
  assign n7570 = n7569 ^ n6356 ;
  assign n7782 = n7635 ^ n7570 ;
  assign n7784 = n7782 ^ x399 ;
  assign n7783 = n7782 ^ n7776 ;
  assign n7785 = n7784 ^ n7783 ;
  assign n7786 = n7781 & ~n7785 ;
  assign n7787 = n7786 ^ n7784 ;
  assign n7914 = n7787 ^ x398 ;
  assign n7915 = ~n7913 & n7914 ;
  assign n7634 = n7633 ^ n7570 ;
  assign n7636 = n7634 & n7635 ;
  assign n7637 = n7636 ^ n5469 ;
  assign n7639 = n7637 ^ n5466 ;
  assign n7365 = ~n7327 & n7364 ;
  assign n7144 = n6434 ^ n5788 ;
  assign n6223 = n6222 ^ n5962 ;
  assign n6848 = n6223 & n6847 ;
  assign n6849 = n6848 ^ n6222 ;
  assign n5961 = n5960 ^ n5955 ;
  assign n6850 = n6849 ^ n5961 ;
  assign n7145 = n6850 ^ n6434 ;
  assign n7146 = ~n7144 & n7145 ;
  assign n7147 = n7146 ^ n5788 ;
  assign n7139 = n7132 ^ n7127 ;
  assign n7140 = n7132 ^ n5021 ;
  assign n7141 = n7139 & n7140 ;
  assign n7142 = n7141 ^ n5021 ;
  assign n7143 = n7142 ^ n5028 ;
  assign n7148 = n7147 ^ n7143 ;
  assign n7150 = n7148 ^ x372 ;
  assign n7149 = n7148 ^ n7133 ;
  assign n7151 = n7150 ^ n7149 ;
  assign n7152 = ~n7138 & n7151 ;
  assign n7153 = n7152 ^ n7150 ;
  assign n7326 = n7153 ^ x371 ;
  assign n7437 = n7365 ^ n7326 ;
  assign n7389 = n7388 ^ n6945 ;
  assign n7433 = n7432 ^ n7388 ;
  assign n7434 = ~n7389 & ~n7433 ;
  assign n7435 = n7434 ^ n6945 ;
  assign n7436 = n7435 ^ n6952 ;
  assign n7564 = n7437 ^ n7436 ;
  assign n7565 = n6805 & n7564 ;
  assign n7566 = n7565 ^ n6364 ;
  assign n7788 = n7639 ^ n7566 ;
  assign n7790 = n7788 ^ x398 ;
  assign n7789 = n7788 ^ n7782 ;
  assign n7791 = n7790 ^ n7789 ;
  assign n7792 = ~n7787 & n7791 ;
  assign n7793 = n7792 ^ n7790 ;
  assign n7916 = n7793 ^ x397 ;
  assign n7917 = n7915 & n7916 ;
  assign n7638 = n7637 ^ n7566 ;
  assign n7640 = ~n7638 & ~n7639 ;
  assign n7641 = n7640 ^ n5466 ;
  assign n7643 = n7641 ^ n5612 ;
  assign n7438 = n7437 ^ n7435 ;
  assign n7439 = n7436 & n7438 ;
  assign n7440 = n7439 ^ n6952 ;
  assign n7560 = n7440 ^ n6877 ;
  assign n7154 = n7147 ^ n7142 ;
  assign n7155 = n6442 ^ n5853 ;
  assign n6856 = n6696 ^ n6695 ;
  assign n6852 = n6442 ^ n6434 ;
  assign n6851 = n6849 ^ n6442 ;
  assign n6853 = n6852 ^ n6851 ;
  assign n6854 = ~n6850 & ~n6853 ;
  assign n6855 = n6854 ^ n6852 ;
  assign n7156 = n6856 ^ n6855 ;
  assign n7157 = n7155 & n7156 ;
  assign n7158 = n7157 ^ n5853 ;
  assign n7159 = n7158 ^ n5028 ;
  assign n7160 = n7159 ^ n7158 ;
  assign n7161 = n7160 ^ n7142 ;
  assign n7162 = ~n7154 & ~n7161 ;
  assign n7163 = n7162 ^ n7159 ;
  assign n7164 = n7163 ^ n5036 ;
  assign n7166 = n7164 ^ x371 ;
  assign n7165 = n7164 ^ n7148 ;
  assign n7167 = n7166 ^ n7165 ;
  assign n7168 = ~n7153 & n7167 ;
  assign n7169 = n7168 ^ n7166 ;
  assign n7367 = n7169 ^ x370 ;
  assign n7366 = ~n7326 & n7365 ;
  assign n7386 = n7367 ^ n7366 ;
  assign n7561 = n7560 ^ n7386 ;
  assign n7562 = n6808 & n7561 ;
  assign n7563 = n7562 ^ n6373 ;
  assign n7794 = n7643 ^ n7563 ;
  assign n7796 = n7794 ^ x397 ;
  assign n7795 = n7794 ^ n7788 ;
  assign n7797 = n7796 ^ n7795 ;
  assign n7798 = ~n7793 & n7797 ;
  assign n7799 = n7798 ^ n7796 ;
  assign n7918 = n7799 ^ x396 ;
  assign n7919 = n7917 & n7918 ;
  assign n7642 = n7641 ^ n7563 ;
  assign n7644 = n7642 & ~n7643 ;
  assign n7645 = n7644 ^ n5612 ;
  assign n7647 = n7645 ^ n5634 ;
  assign n7174 = n6450 ^ n5879 ;
  assign n6862 = n6698 ^ n6697 ;
  assign n6858 = n6450 ^ n6442 ;
  assign n6857 = n6856 ^ n6450 ;
  assign n6859 = n6858 ^ n6857 ;
  assign n6860 = n6855 & n6859 ;
  assign n6861 = n6860 ^ n6858 ;
  assign n7175 = n6862 ^ n6861 ;
  assign n7176 = ~n7174 & ~n7175 ;
  assign n7177 = n7176 ^ n5879 ;
  assign n7170 = n7158 ^ n5036 ;
  assign n7171 = ~n7163 & ~n7170 ;
  assign n7172 = n7171 ^ n5036 ;
  assign n7173 = n7172 ^ n5044 ;
  assign n7178 = n7177 ^ n7173 ;
  assign n7180 = n7178 ^ x370 ;
  assign n7179 = n7178 ^ n7164 ;
  assign n7181 = n7180 ^ n7179 ;
  assign n7182 = n7169 & ~n7181 ;
  assign n7183 = n7182 ^ n7180 ;
  assign n7369 = n7183 ^ x369 ;
  assign n7368 = ~n7366 & ~n7367 ;
  assign n7445 = n7369 ^ n7368 ;
  assign n7387 = n7386 ^ n6877 ;
  assign n7441 = n7440 ^ n7386 ;
  assign n7442 = ~n7387 & n7441 ;
  assign n7443 = n7442 ^ n6877 ;
  assign n7444 = n7443 ^ n6872 ;
  assign n7557 = n7445 ^ n7444 ;
  assign n7558 = n6813 & n7557 ;
  assign n7559 = n7558 ^ n6380 ;
  assign n7800 = n7647 ^ n7559 ;
  assign n7802 = n7800 ^ x396 ;
  assign n7801 = n7800 ^ n7794 ;
  assign n7803 = n7802 ^ n7801 ;
  assign n7804 = ~n7799 & n7803 ;
  assign n7805 = n7804 ^ n7802 ;
  assign n7920 = n7805 ^ x395 ;
  assign n7921 = ~n7919 & ~n7920 ;
  assign n7646 = n7645 ^ n7559 ;
  assign n7648 = n7646 & n7647 ;
  assign n7649 = n7648 ^ n5634 ;
  assign n7651 = n7649 ^ n5650 ;
  assign n7446 = n7445 ^ n7443 ;
  assign n7447 = ~n7444 & ~n7446 ;
  assign n7448 = n7447 ^ n6872 ;
  assign n7553 = n7448 ^ n6967 ;
  assign n7184 = n7177 ^ n7172 ;
  assign n6868 = n6700 ^ n6699 ;
  assign n6864 = n6458 ^ n6450 ;
  assign n6863 = n6862 ^ n6458 ;
  assign n6865 = n6864 ^ n6863 ;
  assign n6866 = n6861 & ~n6865 ;
  assign n6867 = n6866 ^ n6864 ;
  assign n6869 = n6868 ^ n6867 ;
  assign n7185 = n6458 ^ n5907 ;
  assign n7186 = n6869 & ~n7185 ;
  assign n7187 = n7186 ^ n5907 ;
  assign n7188 = n7187 ^ n5044 ;
  assign n7189 = n7188 ^ n7172 ;
  assign n7190 = n7189 ^ n7187 ;
  assign n7191 = ~n7184 & ~n7190 ;
  assign n7192 = n7191 ^ n7188 ;
  assign n7193 = n7192 ^ n5052 ;
  assign n7195 = n7193 ^ x369 ;
  assign n7194 = n7193 ^ n7178 ;
  assign n7196 = n7195 ^ n7194 ;
  assign n7197 = ~n7183 & n7196 ;
  assign n7198 = n7197 ^ n7195 ;
  assign n7371 = n7198 ^ x368 ;
  assign n7370 = ~n7368 & ~n7369 ;
  assign n7384 = n7371 ^ n7370 ;
  assign n7554 = n7553 ^ n7384 ;
  assign n7555 = ~n6817 & ~n7554 ;
  assign n7556 = n7555 ^ n6307 ;
  assign n7806 = n7651 ^ n7556 ;
  assign n7808 = n7806 ^ x395 ;
  assign n7807 = n7806 ^ n7800 ;
  assign n7809 = n7808 ^ n7807 ;
  assign n7810 = ~n7805 & n7809 ;
  assign n7811 = n7810 ^ n7808 ;
  assign n7922 = n7811 ^ x394 ;
  assign n7923 = ~n7921 & n7922 ;
  assign n7650 = n7649 ^ n7556 ;
  assign n7652 = ~n7650 & ~n7651 ;
  assign n7653 = n7652 ^ n5650 ;
  assign n7655 = n7653 ^ n5670 ;
  assign n7199 = n6463 ^ n5973 ;
  assign n7205 = n6702 ^ n6701 ;
  assign n7201 = n6463 ^ n6458 ;
  assign n7200 = n6868 ^ n6463 ;
  assign n7202 = n7201 ^ n7200 ;
  assign n7203 = ~n6867 & n7202 ;
  assign n7204 = n7203 ^ n7201 ;
  assign n7206 = n7205 ^ n7204 ;
  assign n7207 = n7199 & n7206 ;
  assign n7208 = n7207 ^ n5973 ;
  assign n7210 = n7208 ^ n5052 ;
  assign n7209 = n7208 ^ n7187 ;
  assign n7211 = n7210 ^ n7209 ;
  assign n7212 = ~n7192 & n7211 ;
  assign n7213 = n7212 ^ n7210 ;
  assign n7214 = n7213 ^ n4873 ;
  assign n7216 = n7214 ^ x368 ;
  assign n7215 = n7214 ^ n7193 ;
  assign n7217 = n7216 ^ n7215 ;
  assign n7218 = ~n7198 & n7217 ;
  assign n7219 = n7218 ^ n7216 ;
  assign n7373 = n7219 ^ x383 ;
  assign n7372 = ~n7370 & n7371 ;
  assign n7453 = n7373 ^ n7372 ;
  assign n7385 = n7384 ^ n6967 ;
  assign n7449 = n7448 ^ n7384 ;
  assign n7450 = ~n7385 & n7449 ;
  assign n7451 = n7450 ^ n6967 ;
  assign n7452 = n7451 ^ n6977 ;
  assign n7550 = n7453 ^ n7452 ;
  assign n7551 = ~n6822 & n7550 ;
  assign n7552 = n7551 ^ n6392 ;
  assign n7812 = n7655 ^ n7552 ;
  assign n7814 = n7812 ^ x394 ;
  assign n7813 = n7812 ^ n7806 ;
  assign n7815 = n7814 ^ n7813 ;
  assign n7816 = ~n7811 & n7815 ;
  assign n7817 = n7816 ^ n7814 ;
  assign n7924 = n7817 ^ x393 ;
  assign n7925 = n7923 & ~n7924 ;
  assign n7654 = n7653 ^ n7552 ;
  assign n7656 = ~n7654 & ~n7655 ;
  assign n7657 = n7656 ^ n5670 ;
  assign n7818 = n7657 ^ n5690 ;
  assign n7454 = n7453 ^ n7451 ;
  assign n7455 = ~n7452 & n7454 ;
  assign n7456 = n7455 ^ n6977 ;
  assign n7546 = n7456 ^ n7070 ;
  assign n7374 = ~n7372 & ~n7373 ;
  assign n7221 = n7205 ^ n6463 ;
  assign n7222 = ~n7204 & ~n7221 ;
  assign n7223 = n7222 ^ n6463 ;
  assign n7220 = n6704 ^ n6703 ;
  assign n7224 = n7223 ^ n7220 ;
  assign n7225 = n7224 ^ n6267 ;
  assign n7226 = n6266 & n7225 ;
  assign n7227 = n7226 ^ n6267 ;
  assign n7229 = n7227 ^ n4873 ;
  assign n7228 = n7227 ^ n7208 ;
  assign n7230 = n7229 ^ n7228 ;
  assign n7231 = ~n7213 & n7230 ;
  assign n7232 = n7231 ^ n7229 ;
  assign n7233 = n7232 ^ n6014 ;
  assign n7235 = n7233 ^ x383 ;
  assign n7234 = n7233 ^ n7214 ;
  assign n7236 = n7235 ^ n7234 ;
  assign n7237 = ~n7219 & n7236 ;
  assign n7238 = n7237 ^ n7235 ;
  assign n7325 = n7238 ^ x382 ;
  assign n7457 = n7374 ^ n7325 ;
  assign n7547 = n7546 ^ n7457 ;
  assign n7548 = n6828 & n7547 ;
  assign n7549 = n7548 ^ n6399 ;
  assign n7819 = n7818 ^ n7549 ;
  assign n7821 = n7819 ^ x393 ;
  assign n7820 = n7819 ^ n7812 ;
  assign n7822 = n7821 ^ n7820 ;
  assign n7823 = n7817 & ~n7822 ;
  assign n7824 = n7823 ^ n7821 ;
  assign n7926 = n7824 ^ x392 ;
  assign n7927 = n7925 & ~n7926 ;
  assign n7658 = n7657 ^ n7549 ;
  assign n7458 = n7457 ^ n7456 ;
  assign n7459 = n7457 ^ n7070 ;
  assign n7460 = ~n7458 & ~n7459 ;
  assign n7461 = n7460 ^ n7070 ;
  assign n7659 = n7461 ^ n7081 ;
  assign n7375 = n7325 & ~n7374 ;
  assign n7239 = n6298 ^ n6020 ;
  assign n7245 = n6706 ^ n6705 ;
  assign n7243 = n7220 ^ n6298 ;
  assign n7240 = n6267 ^ n6266 ;
  assign n7241 = n7240 ^ n7220 ;
  assign n7242 = ~n7224 & ~n7241 ;
  assign n7244 = n7243 ^ n7242 ;
  assign n7246 = n7245 ^ n7244 ;
  assign n7247 = n7239 & n7246 ;
  assign n7248 = n7247 ^ n6020 ;
  assign n7250 = n7248 ^ n6014 ;
  assign n7249 = n7248 ^ n7227 ;
  assign n7251 = n7250 ^ n7249 ;
  assign n7252 = ~n7232 & n7251 ;
  assign n7253 = n7252 ^ n7250 ;
  assign n7254 = n7253 ^ n5082 ;
  assign n7256 = n7254 ^ x382 ;
  assign n7255 = n7254 ^ n7233 ;
  assign n7257 = n7256 ^ n7255 ;
  assign n7258 = ~n7238 & n7257 ;
  assign n7259 = n7258 ^ n7256 ;
  assign n7324 = n7259 ^ x381 ;
  assign n7462 = n7375 ^ n7324 ;
  assign n7660 = n7659 ^ n7462 ;
  assign n7661 = ~n6833 & n7660 ;
  assign n7662 = n7661 ^ n6407 ;
  assign n7663 = n7662 ^ n5690 ;
  assign n7664 = n7663 ^ n7549 ;
  assign n7665 = n7664 ^ n7662 ;
  assign n7666 = n7658 & n7665 ;
  assign n7667 = n7666 ^ n7663 ;
  assign n7825 = n7667 ^ n5709 ;
  assign n7827 = n7825 ^ x392 ;
  assign n7826 = n7825 ^ n7819 ;
  assign n7828 = n7827 ^ n7826 ;
  assign n7829 = n7824 & ~n7828 ;
  assign n7830 = n7829 ^ n7827 ;
  assign n7928 = n7830 ^ x407 ;
  assign n7929 = n7927 & ~n7928 ;
  assign n7376 = ~n7324 & n7375 ;
  assign n7266 = n6708 ^ n6707 ;
  assign n7260 = n6277 ^ n6276 ;
  assign n7261 = n7260 ^ n6298 ;
  assign n7262 = n7261 ^ n7245 ;
  assign n7263 = n7262 ^ n7260 ;
  assign n7264 = n7244 & ~n7263 ;
  assign n7265 = n7264 ^ n7261 ;
  assign n7267 = n7266 ^ n7265 ;
  assign n7268 = n6276 & ~n7267 ;
  assign n7269 = n7268 ^ n6277 ;
  assign n7271 = n7269 ^ n5082 ;
  assign n7270 = n7269 ^ n7248 ;
  assign n7272 = n7271 ^ n7270 ;
  assign n7273 = n7253 & ~n7272 ;
  assign n7274 = n7273 ^ n7271 ;
  assign n7275 = n7274 ^ n5265 ;
  assign n7277 = n7275 ^ x381 ;
  assign n7276 = n7275 ^ n7254 ;
  assign n7278 = n7277 ^ n7276 ;
  assign n7279 = n7259 & ~n7278 ;
  assign n7280 = n7279 ^ n7277 ;
  assign n7323 = n7280 ^ x380 ;
  assign n7468 = n7376 ^ n7323 ;
  assign n7463 = n7462 ^ n7461 ;
  assign n7464 = n7462 ^ n7081 ;
  assign n7465 = n7463 & n7464 ;
  assign n7466 = n7465 ^ n7081 ;
  assign n7383 = n7095 ^ n6224 ;
  assign n7467 = n7466 ^ n7383 ;
  assign n7542 = n7468 ^ n7467 ;
  assign n7543 = n7095 & ~n7542 ;
  assign n7544 = n7543 ^ n6224 ;
  assign n7669 = n7544 ^ n5709 ;
  assign n7668 = n7662 ^ n7544 ;
  assign n7670 = n7669 ^ n7668 ;
  assign n7671 = ~n7667 & ~n7670 ;
  assign n7672 = n7671 ^ n7669 ;
  assign n7831 = n7672 ^ n5724 ;
  assign n7833 = n7831 ^ x407 ;
  assign n7832 = n7831 ^ n7825 ;
  assign n7834 = n7833 ^ n7832 ;
  assign n7835 = n7830 & ~n7834 ;
  assign n7836 = n7835 ^ n7833 ;
  assign n7930 = n7836 ^ x406 ;
  assign n7931 = n7929 & n7930 ;
  assign n7469 = n7468 ^ n7383 ;
  assign n7470 = n7467 & ~n7469 ;
  assign n7471 = n7470 ^ n7466 ;
  assign n7676 = n7471 ^ n7115 ;
  assign n7377 = ~n7323 & ~n7376 ;
  assign n7285 = n6494 ^ n6064 ;
  assign n7288 = n7266 ^ n7260 ;
  assign n7289 = ~n7265 & n7288 ;
  assign n7287 = n7260 ^ n6494 ;
  assign n7290 = n7289 ^ n7287 ;
  assign n7286 = n6710 ^ n6709 ;
  assign n7291 = n7290 ^ n7286 ;
  assign n7292 = ~n7285 & n7291 ;
  assign n7293 = n7292 ^ n6064 ;
  assign n7281 = n7269 ^ n5265 ;
  assign n7282 = ~n7274 & n7281 ;
  assign n7283 = n7282 ^ n5265 ;
  assign n7284 = n7283 ^ n5286 ;
  assign n7294 = n7293 ^ n7284 ;
  assign n7296 = n7294 ^ x380 ;
  assign n7295 = n7294 ^ n7275 ;
  assign n7297 = n7296 ^ n7295 ;
  assign n7298 = ~n7280 & n7297 ;
  assign n7299 = n7298 ^ n7296 ;
  assign n7322 = n7299 ^ x379 ;
  assign n7381 = n7377 ^ n7322 ;
  assign n7677 = n7676 ^ n7381 ;
  assign n7678 = n6842 & n7677 ;
  assign n7679 = n7678 ^ n6419 ;
  assign n7545 = n7544 ^ n5724 ;
  assign n7673 = ~n7545 & ~n7672 ;
  assign n7674 = n7673 ^ n5724 ;
  assign n7675 = n7674 ^ n5748 ;
  assign n7837 = n7679 ^ n7675 ;
  assign n7839 = n7837 ^ x406 ;
  assign n7838 = n7837 ^ n7831 ;
  assign n7840 = n7839 ^ n7838 ;
  assign n7841 = ~n7836 & n7840 ;
  assign n7842 = n7841 ^ n7839 ;
  assign n7932 = n7842 ^ x405 ;
  assign n7933 = n7931 & n7932 ;
  assign n7684 = n7130 ^ n6222 ;
  assign n7382 = n7381 ^ n7115 ;
  assign n7472 = n7471 ^ n7381 ;
  assign n7473 = ~n7382 & n7472 ;
  assign n7474 = n7473 ^ n7115 ;
  assign n7685 = n7474 ^ n7130 ;
  assign n7378 = ~n7322 & ~n7377 ;
  assign n7305 = n6502 ^ n6117 ;
  assign n7311 = n6712 ^ n6711 ;
  assign n7306 = n6502 ^ n6494 ;
  assign n7307 = n7306 ^ n6502 ;
  assign n7308 = n7307 ^ n7286 ;
  assign n7309 = n7290 & n7308 ;
  assign n7310 = n7309 ^ n7306 ;
  assign n7312 = n7311 ^ n7310 ;
  assign n7313 = ~n7305 & ~n7312 ;
  assign n7314 = n7313 ^ n6117 ;
  assign n7300 = n7293 ^ n7283 ;
  assign n7301 = n7293 ^ n5286 ;
  assign n7302 = n7300 & ~n7301 ;
  assign n7303 = n7302 ^ n5286 ;
  assign n7304 = n7303 ^ n5377 ;
  assign n7315 = n7314 ^ n7304 ;
  assign n7317 = n7315 ^ x379 ;
  assign n7316 = n7315 ^ n7294 ;
  assign n7318 = n7317 ^ n7316 ;
  assign n7319 = n7299 & ~n7318 ;
  assign n7320 = n7319 ^ n7317 ;
  assign n7321 = n7320 ^ x378 ;
  assign n7379 = n7378 ^ n7321 ;
  assign n7686 = n7685 ^ n7379 ;
  assign n7687 = n7684 & ~n7686 ;
  assign n7688 = n7687 ^ n6222 ;
  assign n7680 = n7679 ^ n7674 ;
  assign n7681 = ~n7675 & n7680 ;
  assign n7682 = n7681 ^ n5748 ;
  assign n7683 = n7682 ^ n5768 ;
  assign n7843 = n7688 ^ n7683 ;
  assign n7845 = n7843 ^ x405 ;
  assign n7844 = n7843 ^ n7837 ;
  assign n7846 = n7845 ^ n7844 ;
  assign n7847 = ~n7842 & n7846 ;
  assign n7848 = n7847 ^ n7845 ;
  assign n7934 = n7848 ^ x404 ;
  assign n7935 = n7933 & ~n7934 ;
  assign n7380 = n7379 ^ n7130 ;
  assign n7475 = n7474 ^ n7379 ;
  assign n7476 = n7380 & ~n7475 ;
  assign n7477 = n7476 ^ n7130 ;
  assign n7693 = n7477 ^ n7145 ;
  assign n7500 = ~n7321 & n7378 ;
  assign n7483 = n6510 ^ n6143 ;
  assign n7489 = n6714 ^ n6713 ;
  assign n7485 = n6510 ^ n6502 ;
  assign n7484 = n7311 ^ n6510 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7487 = ~n7310 & ~n7486 ;
  assign n7488 = n7487 ^ n7485 ;
  assign n7490 = n7489 ^ n7488 ;
  assign n7491 = n7483 & ~n7490 ;
  assign n7492 = n7491 ^ n6143 ;
  assign n7478 = n7314 ^ n7303 ;
  assign n7479 = n7314 ^ n5377 ;
  assign n7480 = ~n7478 & ~n7479 ;
  assign n7481 = n7480 ^ n5377 ;
  assign n7482 = n7481 ^ n5408 ;
  assign n7493 = n7492 ^ n7482 ;
  assign n7495 = n7493 ^ x378 ;
  assign n7494 = n7493 ^ n7315 ;
  assign n7496 = n7495 ^ n7494 ;
  assign n7497 = n7320 & ~n7496 ;
  assign n7498 = n7497 ^ n7495 ;
  assign n7499 = n7498 ^ x377 ;
  assign n7501 = n7500 ^ n7499 ;
  assign n7694 = n7693 ^ n7501 ;
  assign n7695 = n6850 & ~n7694 ;
  assign n7696 = n7695 ^ n6434 ;
  assign n7689 = n7688 ^ n7682 ;
  assign n7690 = n7683 & ~n7689 ;
  assign n7691 = n7690 ^ n5768 ;
  assign n7692 = n7691 ^ n5788 ;
  assign n7849 = n7696 ^ n7692 ;
  assign n7851 = n7849 ^ x404 ;
  assign n7850 = n7849 ^ n7843 ;
  assign n7852 = n7851 ^ n7850 ;
  assign n7853 = n7848 & ~n7852 ;
  assign n7854 = n7853 ^ n7851 ;
  assign n7936 = n7854 ^ x403 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7701 = n7156 ^ n6442 ;
  assign n7502 = n7501 ^ n7477 ;
  assign n7503 = n7501 ^ n7145 ;
  assign n7504 = n7502 & n7503 ;
  assign n7505 = n7504 ^ n7145 ;
  assign n7702 = n7505 ^ n7156 ;
  assign n7523 = n7500 ^ n7493 ;
  assign n7524 = ~n7498 & ~n7523 ;
  assign n7521 = n7500 ^ n7498 ;
  assign n7522 = ~x377 & n7521 ;
  assign n7525 = n7524 ^ n7522 ;
  assign n7517 = n5408 ^ x376 ;
  assign n7518 = n7517 ^ n6225 ;
  assign n7509 = n6295 ^ n6171 ;
  assign n7513 = n7489 ^ n6510 ;
  assign n7514 = n7488 & n7513 ;
  assign n7511 = n6716 ^ n6715 ;
  assign n7510 = n7489 ^ n6295 ;
  assign n7512 = n7511 ^ n7510 ;
  assign n7515 = n7514 ^ n7512 ;
  assign n7516 = ~n7509 & ~n7515 ;
  assign n7519 = n7518 ^ n7516 ;
  assign n7506 = n7492 ^ n7481 ;
  assign n7507 = n7492 ^ n5408 ;
  assign n7508 = n7506 & ~n7507 ;
  assign n7520 = n7519 ^ n7508 ;
  assign n7526 = n7525 ^ n7520 ;
  assign n7703 = n7702 ^ n7526 ;
  assign n7704 = n7701 & n7703 ;
  assign n7705 = n7704 ^ n6442 ;
  assign n7697 = n7696 ^ n7691 ;
  assign n7698 = n7692 & n7697 ;
  assign n7699 = n7698 ^ n5788 ;
  assign n7700 = n7699 ^ n5853 ;
  assign n7855 = n7705 ^ n7700 ;
  assign n7857 = n7855 ^ x403 ;
  assign n7856 = n7855 ^ n7849 ;
  assign n7858 = n7857 ^ n7856 ;
  assign n7859 = ~n7854 & n7858 ;
  assign n7860 = n7859 ^ n7857 ;
  assign n7938 = n7860 ^ x402 ;
  assign n7939 = ~n7937 & ~n7938 ;
  assign n7710 = n7175 ^ n6450 ;
  assign n7533 = n6985 ^ x359 ;
  assign n7527 = n7526 ^ n7505 ;
  assign n7528 = n7175 ^ n7156 ;
  assign n7529 = n7528 ^ n7175 ;
  assign n7530 = n7529 ^ n7505 ;
  assign n7531 = ~n7527 & n7530 ;
  assign n7532 = n7531 ^ n7528 ;
  assign n7711 = n7533 ^ n7532 ;
  assign n7712 = ~n7710 & n7711 ;
  assign n7713 = n7712 ^ n6450 ;
  assign n7706 = n7705 ^ n7699 ;
  assign n7707 = ~n7700 & n7706 ;
  assign n7708 = n7707 ^ n5853 ;
  assign n7709 = n7708 ^ n5879 ;
  assign n7861 = n7713 ^ n7709 ;
  assign n7863 = n7861 ^ x402 ;
  assign n7862 = n7861 ^ n7855 ;
  assign n7864 = n7863 ^ n7862 ;
  assign n7865 = n7860 & ~n7864 ;
  assign n7866 = n7865 ^ n7863 ;
  assign n7940 = n7866 ^ x401 ;
  assign n7941 = n7939 & ~n7940 ;
  assign n7714 = n7713 ^ n7708 ;
  assign n7715 = ~n7709 & ~n7714 ;
  assign n7716 = n7715 ^ n5879 ;
  assign n7733 = n7716 ^ n5907 ;
  assign n6870 = n6869 ^ n6458 ;
  assign n7535 = n7175 ^ n6869 ;
  assign n7534 = n7533 ^ n6869 ;
  assign n7536 = n7535 ^ n7534 ;
  assign n7537 = ~n7532 & n7536 ;
  assign n7538 = n7537 ^ n7535 ;
  assign n7539 = n7538 ^ n7332 ;
  assign n7540 = ~n6870 & n7539 ;
  assign n7541 = n7540 ^ n6458 ;
  assign n7734 = n7733 ^ n7541 ;
  assign n7868 = n7734 ^ x401 ;
  assign n7867 = n7861 ^ n7734 ;
  assign n7869 = n7868 ^ n7867 ;
  assign n7870 = n7866 & ~n7869 ;
  assign n7871 = n7870 ^ n7868 ;
  assign n7942 = n7871 ^ x400 ;
  assign n7943 = ~n7941 & ~n7942 ;
  assign n7735 = n7734 ^ x400 ;
  assign n7872 = n7735 & ~n7871 ;
  assign n7873 = n7872 ^ x400 ;
  assign n7717 = n7716 ^ n7541 ;
  assign n7718 = n7206 ^ n6463 ;
  assign n7722 = n7333 ^ n7332 ;
  assign n7723 = n7722 ^ n7206 ;
  assign n7719 = n7332 ^ n6869 ;
  assign n7720 = n7538 & ~n7719 ;
  assign n7721 = n7720 ^ n7332 ;
  assign n7724 = n7723 ^ n7721 ;
  assign n7725 = n7718 & ~n7724 ;
  assign n7726 = n7725 ^ n6463 ;
  assign n7727 = n7726 ^ n5907 ;
  assign n7728 = n7727 ^ n7541 ;
  assign n7729 = n7728 ^ n7726 ;
  assign n7730 = ~n7717 & ~n7729 ;
  assign n7731 = n7730 ^ n7727 ;
  assign n7732 = n7731 ^ n5973 ;
  assign n7874 = n7873 ^ n7732 ;
  assign n7944 = n7874 ^ x415 ;
  assign n7945 = n7943 & ~n7944 ;
  assign n7882 = n7335 ^ n7334 ;
  assign n7875 = n7722 ^ n7721 ;
  assign n7876 = n7240 ^ n7224 ;
  assign n7877 = n7876 ^ n7206 ;
  assign n7878 = n7877 ^ n7721 ;
  assign n7879 = n7878 ^ n7876 ;
  assign n7880 = n7875 & ~n7879 ;
  assign n7881 = n7880 ^ n7877 ;
  assign n7883 = n7882 ^ n7881 ;
  assign n7884 = ~n7224 & n7883 ;
  assign n7885 = n7884 ^ n7240 ;
  assign n7887 = n7885 ^ n5973 ;
  assign n7886 = n7885 ^ n7726 ;
  assign n7888 = n7887 ^ n7886 ;
  assign n7889 = ~n7731 & n7888 ;
  assign n7890 = n7889 ^ n7887 ;
  assign n7891 = n7890 ^ n6267 ;
  assign n7892 = n7891 ^ x415 ;
  assign n7893 = n7892 ^ n7873 ;
  assign n7894 = n7893 ^ n7891 ;
  assign n7895 = ~n7874 & n7894 ;
  assign n7896 = n7895 ^ n7892 ;
  assign n7897 = n7896 ^ x414 ;
  assign n7946 = n7945 ^ n7897 ;
  assign n8520 = n7974 ^ n7946 ;
  assign n7947 = n7946 ^ n7395 ;
  assign n7948 = ~n7396 & n7947 ;
  assign n7949 = n7948 ^ n7395 ;
  assign n7981 = n7949 ^ n6763 ;
  assign n7982 = x423 & ~n7981 ;
  assign n7975 = n7946 & n7974 ;
  assign n7976 = n7975 ^ n7595 ;
  assign n7972 = ~n7897 & n7945 ;
  assign n7956 = n7246 ^ n6298 ;
  assign n7959 = n7882 ^ n7876 ;
  assign n7960 = ~n7881 & n7959 ;
  assign n7958 = n7876 ^ n7246 ;
  assign n7961 = n7960 ^ n7958 ;
  assign n7957 = n7337 ^ n7336 ;
  assign n7962 = n7961 ^ n7957 ;
  assign n7963 = ~n7956 & ~n7962 ;
  assign n7964 = n7963 ^ n6298 ;
  assign n7952 = n7885 ^ n6267 ;
  assign n7953 = ~n7890 & n7952 ;
  assign n7954 = n7953 ^ n6267 ;
  assign n7955 = n7954 ^ n6020 ;
  assign n7965 = n7964 ^ n7955 ;
  assign n7967 = n7965 ^ x414 ;
  assign n7966 = n7965 ^ n7891 ;
  assign n7968 = n7967 ^ n7966 ;
  assign n7969 = ~n7896 & n7968 ;
  assign n7970 = n7969 ^ n7967 ;
  assign n7971 = n7970 ^ x413 ;
  assign n7973 = n7972 ^ n7971 ;
  assign n7977 = n7976 ^ n7973 ;
  assign n7978 = ~n7400 & ~n7977 ;
  assign n7979 = n7978 ^ n6885 ;
  assign n7950 = n6763 & ~n7949 ;
  assign n7951 = n7950 ^ n5927 ;
  assign n7980 = n7979 ^ n7951 ;
  assign n7983 = n7982 ^ n7980 ;
  assign n8012 = n7975 ^ n7973 ;
  assign n8013 = n7976 & n8012 ;
  assign n8014 = n8013 ^ n7595 ;
  assign n8015 = n8014 ^ n7592 ;
  assign n8010 = n7971 & ~n7972 ;
  assign n7993 = n7267 ^ n7260 ;
  assign n7999 = n7339 ^ n7338 ;
  assign n7994 = n7267 ^ n7246 ;
  assign n7995 = n7994 ^ n7267 ;
  assign n7996 = n7995 ^ n7957 ;
  assign n7997 = ~n7961 & n7996 ;
  assign n7998 = n7997 ^ n7994 ;
  assign n8000 = n7999 ^ n7998 ;
  assign n8001 = ~n7993 & ~n8000 ;
  assign n8002 = n8001 ^ n7260 ;
  assign n7988 = n7964 ^ n7954 ;
  assign n7989 = n7964 ^ n6020 ;
  assign n7990 = n7988 & n7989 ;
  assign n7991 = n7990 ^ n6020 ;
  assign n7992 = n7991 ^ n6277 ;
  assign n8003 = n8002 ^ n7992 ;
  assign n8005 = n8003 ^ x413 ;
  assign n8004 = n8003 ^ n7965 ;
  assign n8006 = n8005 ^ n8004 ;
  assign n8007 = ~n7970 & n8006 ;
  assign n8008 = n8007 ^ n8005 ;
  assign n8009 = n8008 ^ x412 ;
  assign n8011 = n8010 ^ n8009 ;
  assign n8016 = n8015 ^ n8011 ;
  assign n8017 = n7405 & n8016 ;
  assign n8018 = n8017 ^ n6892 ;
  assign n7984 = n7979 ^ n7950 ;
  assign n7985 = n7951 & n7984 ;
  assign n7986 = n7985 ^ n5927 ;
  assign n7987 = n7986 ^ n5934 ;
  assign n8019 = n8018 ^ n7987 ;
  assign n8020 = n8019 ^ x422 ;
  assign n8021 = n8020 ^ n7980 ;
  assign n8022 = n8021 ^ n8019 ;
  assign n8023 = n7983 & ~n8022 ;
  assign n8024 = n8023 ^ n8020 ;
  assign n8061 = n8009 & ~n8010 ;
  assign n8044 = n7291 ^ n6494 ;
  assign n8050 = n7341 ^ n7340 ;
  assign n8046 = n7291 ^ n7267 ;
  assign n8045 = n7999 ^ n7291 ;
  assign n8047 = n8046 ^ n8045 ;
  assign n8048 = ~n7998 & ~n8047 ;
  assign n8049 = n8048 ^ n8046 ;
  assign n8051 = n8050 ^ n8049 ;
  assign n8052 = n8044 & n8051 ;
  assign n8053 = n8052 ^ n6494 ;
  assign n8039 = n8002 ^ n7991 ;
  assign n8040 = n8002 ^ n6277 ;
  assign n8041 = n8039 & n8040 ;
  assign n8042 = n8041 ^ n6277 ;
  assign n8043 = n8042 ^ n6064 ;
  assign n8054 = n8053 ^ n8043 ;
  assign n8056 = n8054 ^ x412 ;
  assign n8055 = n8054 ^ n8003 ;
  assign n8057 = n8056 ^ n8055 ;
  assign n8058 = n8008 & ~n8057 ;
  assign n8059 = n8058 ^ n8056 ;
  assign n8060 = n8059 ^ x411 ;
  assign n8062 = n8061 ^ n8060 ;
  assign n8035 = n8014 ^ n8011 ;
  assign n8036 = n8015 & ~n8035 ;
  assign n8037 = n8036 ^ n7592 ;
  assign n8038 = n8037 ^ n7589 ;
  assign n8063 = n8062 ^ n8038 ;
  assign n8064 = n7408 & ~n8063 ;
  assign n8065 = n8064 ^ n6900 ;
  assign n8031 = n8018 ^ n7986 ;
  assign n8032 = ~n7987 & ~n8031 ;
  assign n8033 = n8032 ^ n5934 ;
  assign n8034 = n8033 ^ n5919 ;
  assign n8066 = n8065 ^ n8034 ;
  assign n8068 = n8066 ^ x421 ;
  assign n8067 = n8066 ^ n8019 ;
  assign n8069 = n8068 ^ n8067 ;
  assign n8070 = n8024 & ~n8069 ;
  assign n8071 = n8070 ^ n8068 ;
  assign n8102 = n8062 ^ n7589 ;
  assign n8103 = n8062 ^ n8037 ;
  assign n8104 = ~n8102 & ~n8103 ;
  assign n8105 = n8104 ^ n7589 ;
  assign n8106 = n8105 ^ n7585 ;
  assign n8100 = ~n8060 & ~n8061 ;
  assign n8083 = n7312 ^ n6502 ;
  assign n8089 = n7343 ^ n7342 ;
  assign n8085 = n7312 ^ n7291 ;
  assign n8084 = n8050 ^ n7312 ;
  assign n8086 = n8085 ^ n8084 ;
  assign n8087 = ~n8049 & ~n8086 ;
  assign n8088 = n8087 ^ n8085 ;
  assign n8090 = n8089 ^ n8088 ;
  assign n8091 = n8083 & n8090 ;
  assign n8092 = n8091 ^ n6502 ;
  assign n8078 = n8053 ^ n8042 ;
  assign n8079 = n8053 ^ n6064 ;
  assign n8080 = ~n8078 & ~n8079 ;
  assign n8081 = n8080 ^ n6064 ;
  assign n8082 = n8081 ^ n6117 ;
  assign n8093 = n8092 ^ n8082 ;
  assign n8095 = n8093 ^ x411 ;
  assign n8094 = n8093 ^ n8054 ;
  assign n8096 = n8095 ^ n8094 ;
  assign n8097 = n8059 & ~n8096 ;
  assign n8098 = n8097 ^ n8095 ;
  assign n8099 = n8098 ^ x410 ;
  assign n8101 = n8100 ^ n8099 ;
  assign n8107 = n8106 ^ n8101 ;
  assign n8108 = n7413 & ~n8107 ;
  assign n8109 = n8108 ^ n6907 ;
  assign n8074 = n8065 ^ n8033 ;
  assign n8075 = ~n8034 & ~n8074 ;
  assign n8076 = n8075 ^ n5919 ;
  assign n8077 = n8076 ^ n6315 ;
  assign n8110 = n8109 ^ n8077 ;
  assign n8112 = n8110 ^ x420 ;
  assign n8111 = n8110 ^ n8066 ;
  assign n8113 = n8112 ^ n8111 ;
  assign n8114 = ~n8071 & n8113 ;
  assign n8115 = n8114 ^ n8112 ;
  assign n8132 = n7490 ^ n6510 ;
  assign n8138 = n7345 ^ n7344 ;
  assign n8134 = n7490 ^ n7312 ;
  assign n8133 = n8089 ^ n7490 ;
  assign n8135 = n8134 ^ n8133 ;
  assign n8136 = ~n8088 & n8135 ;
  assign n8137 = n8136 ^ n8134 ;
  assign n8139 = n8138 ^ n8137 ;
  assign n8140 = ~n8132 & n8139 ;
  assign n8141 = n8140 ^ n6510 ;
  assign n8127 = n8092 ^ n8081 ;
  assign n8128 = n8092 ^ n6117 ;
  assign n8129 = ~n8127 & ~n8128 ;
  assign n8130 = n8129 ^ n6117 ;
  assign n8131 = n8130 ^ n6143 ;
  assign n8142 = n8141 ^ n8131 ;
  assign n8144 = n8142 ^ x410 ;
  assign n8143 = n8142 ^ n8093 ;
  assign n8145 = n8144 ^ n8143 ;
  assign n8146 = ~n8098 & n8145 ;
  assign n8147 = n8146 ^ n8144 ;
  assign n8148 = n8147 ^ x409 ;
  assign n8126 = ~n8099 & ~n8100 ;
  assign n8149 = n8148 ^ n8126 ;
  assign n8122 = n8105 ^ n8101 ;
  assign n8123 = n8106 & ~n8122 ;
  assign n8124 = n8123 ^ n7585 ;
  assign n8125 = n8124 ^ n7582 ;
  assign n8150 = n8149 ^ n8125 ;
  assign n8151 = ~n7416 & n8150 ;
  assign n8152 = n8151 ^ n6915 ;
  assign n8118 = n8109 ^ n8076 ;
  assign n8119 = ~n8077 & n8118 ;
  assign n8120 = n8119 ^ n6315 ;
  assign n8121 = n8120 ^ n6322 ;
  assign n8153 = n8152 ^ n8121 ;
  assign n8155 = n8153 ^ x419 ;
  assign n8154 = n8153 ^ n8110 ;
  assign n8156 = n8155 ^ n8154 ;
  assign n8157 = ~n8115 & n8156 ;
  assign n8158 = n8157 ^ n8155 ;
  assign n8181 = n7515 ^ n6295 ;
  assign n8185 = n8138 ^ n7490 ;
  assign n8186 = ~n8137 & ~n8185 ;
  assign n8182 = n7347 ^ n7346 ;
  assign n8183 = n8182 ^ n7515 ;
  assign n8184 = n8183 ^ n8138 ;
  assign n8187 = n8186 ^ n8184 ;
  assign n8188 = ~n8181 & n8187 ;
  assign n8178 = n6143 ^ x408 ;
  assign n8179 = n8178 ^ n7509 ;
  assign n8175 = n8141 ^ n8130 ;
  assign n8176 = n8141 ^ n6143 ;
  assign n8177 = ~n8175 & n8176 ;
  assign n8180 = n8179 ^ n8177 ;
  assign n8189 = n8188 ^ n8180 ;
  assign n8170 = n8142 ^ n8126 ;
  assign n8173 = ~n8147 & n8170 ;
  assign n8169 = n8147 ^ n8142 ;
  assign n8171 = n8170 ^ n8169 ;
  assign n8172 = x409 & n8171 ;
  assign n8174 = n8173 ^ n8172 ;
  assign n8190 = n8189 ^ n8174 ;
  assign n8191 = n8190 ^ n7578 ;
  assign n8165 = n8149 ^ n8124 ;
  assign n8166 = n8149 ^ n7582 ;
  assign n8167 = n8165 & ~n8166 ;
  assign n8168 = n8167 ^ n7582 ;
  assign n8192 = n8191 ^ n8168 ;
  assign n8193 = n7421 & n8192 ;
  assign n8194 = n8193 ^ n6922 ;
  assign n8161 = n8152 ^ n8120 ;
  assign n8162 = n8121 & n8161 ;
  assign n8163 = n8162 ^ n6322 ;
  assign n8164 = n8163 ^ n6330 ;
  assign n8195 = n8194 ^ n8164 ;
  assign n8197 = n8195 ^ x418 ;
  assign n8196 = n8195 ^ n8153 ;
  assign n8198 = n8197 ^ n8196 ;
  assign n8199 = ~n8158 & n8198 ;
  assign n8200 = n8199 ^ n8197 ;
  assign n8214 = n7737 ^ x391 ;
  assign n8208 = n8190 ^ n8168 ;
  assign n8211 = n8168 ^ n7578 ;
  assign n8212 = n8208 & n8211 ;
  assign n8209 = n7578 ^ n7575 ;
  assign n8213 = n8212 ^ n8209 ;
  assign n8215 = n8214 ^ n8213 ;
  assign n8216 = n7424 & n8215 ;
  assign n8217 = n8216 ^ n6930 ;
  assign n8203 = n8194 ^ n6330 ;
  assign n8204 = n8194 ^ n8163 ;
  assign n8205 = ~n8203 & ~n8204 ;
  assign n8206 = n8205 ^ n6330 ;
  assign n8207 = n8206 ^ n6339 ;
  assign n8218 = n8217 ^ n8207 ;
  assign n8220 = n8218 ^ x417 ;
  assign n8219 = n8218 ^ n8195 ;
  assign n8221 = n8220 ^ n8219 ;
  assign n8222 = ~n8200 & n8221 ;
  assign n8223 = n8222 ^ n8220 ;
  assign n8240 = n8218 ^ x416 ;
  assign n8241 = ~n8223 & n8240 ;
  assign n8242 = n8241 ^ x416 ;
  assign n8231 = n8214 ^ n7575 ;
  assign n8232 = n8213 & ~n8231 ;
  assign n8233 = n8232 ^ n7575 ;
  assign n8234 = n8233 ^ n7572 ;
  assign n8235 = n8234 ^ n7900 ;
  assign n8236 = n7429 & ~n8235 ;
  assign n8237 = n8236 ^ n6937 ;
  assign n8226 = n8217 ^ n8206 ;
  assign n8227 = n8217 ^ n6339 ;
  assign n8228 = n8226 & n8227 ;
  assign n8229 = n8228 ^ n6339 ;
  assign n8230 = n8229 ^ n6348 ;
  assign n8238 = n8237 ^ n8230 ;
  assign n8245 = n8242 ^ n8238 ;
  assign n8257 = n7901 ^ n7900 ;
  assign n8251 = n8233 ^ n7900 ;
  assign n8255 = ~n8234 & n8251 ;
  assign n8252 = n7572 ^ n7568 ;
  assign n8256 = n8255 ^ n8252 ;
  assign n8258 = n8257 ^ n8256 ;
  assign n8259 = n7433 & n8258 ;
  assign n8260 = n8259 ^ n6945 ;
  assign n8246 = n8237 ^ n8229 ;
  assign n8247 = n8237 ^ n6348 ;
  assign n8248 = n8246 & ~n8247 ;
  assign n8249 = n8248 ^ n6348 ;
  assign n8250 = n8249 ^ n6356 ;
  assign n8261 = n8260 ^ n8250 ;
  assign n8262 = n8261 ^ x431 ;
  assign n8263 = n8262 ^ n8238 ;
  assign n8264 = n8263 ^ n8261 ;
  assign n8265 = ~n8245 & n8264 ;
  assign n8266 = n8265 ^ n8262 ;
  assign n8279 = n7902 ^ n7898 ;
  assign n8275 = n7568 ^ n7564 ;
  assign n8274 = n8257 ^ n7564 ;
  assign n8276 = n8275 ^ n8274 ;
  assign n8277 = ~n8256 & n8276 ;
  assign n8278 = n8277 ^ n8275 ;
  assign n8280 = n8279 ^ n8278 ;
  assign n8281 = ~n7438 & n8280 ;
  assign n8282 = n8281 ^ n6952 ;
  assign n8269 = n8260 ^ n8249 ;
  assign n8270 = n8260 ^ n6356 ;
  assign n8271 = ~n8269 & ~n8270 ;
  assign n8272 = n8271 ^ n6356 ;
  assign n8273 = n8272 ^ n6364 ;
  assign n8283 = n8282 ^ n8273 ;
  assign n8285 = n8283 ^ x430 ;
  assign n8284 = n8283 ^ n8261 ;
  assign n8286 = n8285 ^ n8284 ;
  assign n8287 = ~n8266 & n8286 ;
  assign n8288 = n8287 ^ n8285 ;
  assign n8291 = n8282 ^ n8272 ;
  assign n8292 = n7904 ^ n7903 ;
  assign n8294 = n8292 ^ n7564 ;
  assign n8293 = n8292 ^ n8279 ;
  assign n8295 = n8294 ^ n8293 ;
  assign n8296 = ~n8278 & ~n8295 ;
  assign n8297 = n8296 ^ n8294 ;
  assign n8298 = n8297 ^ n7561 ;
  assign n8299 = ~n7441 & ~n8298 ;
  assign n8300 = n8299 ^ n6877 ;
  assign n8301 = n8300 ^ n6364 ;
  assign n8302 = n8301 ^ n8300 ;
  assign n8303 = n8302 ^ n8272 ;
  assign n8304 = n8291 & ~n8303 ;
  assign n8305 = n8304 ^ n8301 ;
  assign n8306 = n8305 ^ n6373 ;
  assign n8308 = n8306 ^ x429 ;
  assign n8307 = n8306 ^ n8283 ;
  assign n8309 = n8308 ^ n8307 ;
  assign n8310 = ~n8288 & n8309 ;
  assign n8311 = n8310 ^ n8308 ;
  assign n8323 = n7906 ^ n7905 ;
  assign n8319 = n7561 ^ n7557 ;
  assign n8318 = n8292 ^ n7557 ;
  assign n8320 = n8319 ^ n8318 ;
  assign n8321 = n8297 & ~n8320 ;
  assign n8322 = n8321 ^ n8319 ;
  assign n8324 = n8323 ^ n8322 ;
  assign n8325 = n7446 & ~n8324 ;
  assign n8326 = n8325 ^ n6872 ;
  assign n8314 = n8300 ^ n6373 ;
  assign n8315 = ~n8305 & n8314 ;
  assign n8316 = n8315 ^ n6373 ;
  assign n8317 = n8316 ^ n6380 ;
  assign n8327 = n8326 ^ n8317 ;
  assign n8329 = n8327 ^ x428 ;
  assign n8328 = n8327 ^ n8306 ;
  assign n8330 = n8329 ^ n8328 ;
  assign n8331 = n8311 & ~n8330 ;
  assign n8332 = n8331 ^ n8329 ;
  assign n8345 = n7908 ^ n7907 ;
  assign n8341 = n7557 ^ n7554 ;
  assign n8340 = n8323 ^ n7554 ;
  assign n8342 = n8341 ^ n8340 ;
  assign n8343 = n8322 & ~n8342 ;
  assign n8344 = n8343 ^ n8341 ;
  assign n8346 = n8345 ^ n8344 ;
  assign n8347 = ~n7449 & n8346 ;
  assign n8348 = n8347 ^ n6967 ;
  assign n8335 = n8326 ^ n8316 ;
  assign n8336 = n8326 ^ n6380 ;
  assign n8337 = n8335 & n8336 ;
  assign n8338 = n8337 ^ n6380 ;
  assign n8339 = n8338 ^ n6307 ;
  assign n8349 = n8348 ^ n8339 ;
  assign n8351 = n8349 ^ x427 ;
  assign n8350 = n8349 ^ n8327 ;
  assign n8352 = n8351 ^ n8350 ;
  assign n8353 = n8332 & ~n8352 ;
  assign n8354 = n8353 ^ n8351 ;
  assign n8357 = n8348 ^ n8338 ;
  assign n8363 = n7910 ^ n7909 ;
  assign n8359 = n7554 ^ n7550 ;
  assign n8358 = n8345 ^ n7550 ;
  assign n8360 = n8359 ^ n8358 ;
  assign n8361 = ~n8344 & n8360 ;
  assign n8362 = n8361 ^ n8359 ;
  assign n8364 = n8363 ^ n8362 ;
  assign n8365 = ~n7454 & ~n8364 ;
  assign n8366 = n8365 ^ n6977 ;
  assign n8367 = n8366 ^ n6307 ;
  assign n8368 = n8367 ^ n8366 ;
  assign n8369 = n8368 ^ n8338 ;
  assign n8370 = ~n8357 & ~n8369 ;
  assign n8371 = n8370 ^ n8367 ;
  assign n8372 = n8371 ^ n6392 ;
  assign n8374 = n8372 ^ x426 ;
  assign n8373 = n8372 ^ n8349 ;
  assign n8375 = n8374 ^ n8373 ;
  assign n8376 = n8354 & ~n8375 ;
  assign n8377 = n8376 ^ n8374 ;
  assign n8389 = n7912 ^ n7911 ;
  assign n8385 = n7550 ^ n7547 ;
  assign n8384 = n8363 ^ n7547 ;
  assign n8386 = n8385 ^ n8384 ;
  assign n8387 = ~n8362 & n8386 ;
  assign n8388 = n8387 ^ n8385 ;
  assign n8390 = n8389 ^ n8388 ;
  assign n8391 = n7458 & n8390 ;
  assign n8392 = n8391 ^ n7070 ;
  assign n8380 = n8366 ^ n6392 ;
  assign n8381 = ~n8371 & ~n8380 ;
  assign n8382 = n8381 ^ n6392 ;
  assign n8383 = n8382 ^ n6399 ;
  assign n8393 = n8392 ^ n8383 ;
  assign n8395 = n8393 ^ x425 ;
  assign n8394 = n8393 ^ n8372 ;
  assign n8396 = n8395 ^ n8394 ;
  assign n8397 = ~n8377 & n8396 ;
  assign n8398 = n8397 ^ n8395 ;
  assign n8401 = n8392 ^ n8382 ;
  assign n8407 = n7914 ^ n7913 ;
  assign n8403 = n7660 ^ n7547 ;
  assign n8402 = n8389 ^ n7660 ;
  assign n8404 = n8403 ^ n8402 ;
  assign n8405 = n8388 & n8404 ;
  assign n8406 = n8405 ^ n8403 ;
  assign n8408 = n8407 ^ n8406 ;
  assign n8409 = ~n7463 & ~n8408 ;
  assign n8410 = n8409 ^ n7081 ;
  assign n8411 = n8410 ^ n6399 ;
  assign n8412 = n8411 ^ n8382 ;
  assign n8413 = n8412 ^ n8410 ;
  assign n8414 = ~n8401 & n8413 ;
  assign n8415 = n8414 ^ n8411 ;
  assign n8416 = n8415 ^ n6407 ;
  assign n8418 = n8416 ^ x424 ;
  assign n8417 = n8416 ^ n8393 ;
  assign n8419 = n8418 ^ n8417 ;
  assign n8420 = ~n8398 & n8419 ;
  assign n8421 = n8420 ^ n8418 ;
  assign n8428 = n7468 ^ n7466 ;
  assign n8429 = n7916 ^ n7915 ;
  assign n8431 = n8429 ^ n7660 ;
  assign n8430 = n8429 ^ n8407 ;
  assign n8432 = n8431 ^ n8430 ;
  assign n8433 = n8406 & ~n8432 ;
  assign n8434 = n8433 ^ n8431 ;
  assign n8435 = n8434 ^ n7383 ;
  assign n8436 = n8428 & n8435 ;
  assign n8437 = n8436 ^ n7383 ;
  assign n8424 = n8410 ^ n6407 ;
  assign n8425 = n8415 & ~n8424 ;
  assign n8426 = n8425 ^ n6407 ;
  assign n8427 = n8426 ^ n6224 ;
  assign n8438 = n8437 ^ n8427 ;
  assign n8440 = n8438 ^ x439 ;
  assign n8439 = n8438 ^ n8416 ;
  assign n8441 = n8440 ^ n8439 ;
  assign n8442 = n8421 & ~n8441 ;
  assign n8443 = n8442 ^ n8440 ;
  assign n8446 = n8437 ^ n8426 ;
  assign n8452 = n7918 ^ n7917 ;
  assign n8448 = n7677 ^ n7542 ;
  assign n8447 = n8429 ^ n7677 ;
  assign n8449 = n8448 ^ n8447 ;
  assign n8450 = ~n8434 & ~n8449 ;
  assign n8451 = n8450 ^ n8448 ;
  assign n8453 = n8452 ^ n8451 ;
  assign n8454 = ~n7472 & ~n8453 ;
  assign n8455 = n8454 ^ n7115 ;
  assign n8456 = n8455 ^ n6224 ;
  assign n8457 = n8456 ^ n8426 ;
  assign n8458 = n8457 ^ n8455 ;
  assign n8459 = n8446 & ~n8458 ;
  assign n8460 = n8459 ^ n8456 ;
  assign n8461 = n8460 ^ n6419 ;
  assign n8463 = n8461 ^ x438 ;
  assign n8462 = n8461 ^ n8438 ;
  assign n8464 = n8463 ^ n8462 ;
  assign n8465 = ~n8443 & n8464 ;
  assign n8466 = n8465 ^ n8463 ;
  assign n8478 = n7920 ^ n7919 ;
  assign n8474 = n7686 ^ n7677 ;
  assign n8473 = n8452 ^ n7686 ;
  assign n8475 = n8474 ^ n8473 ;
  assign n8476 = ~n8451 & n8475 ;
  assign n8477 = n8476 ^ n8474 ;
  assign n8479 = n8478 ^ n8477 ;
  assign n8480 = n7475 & n8479 ;
  assign n8481 = n8480 ^ n7130 ;
  assign n8469 = n8455 ^ n6419 ;
  assign n8470 = ~n8460 & n8469 ;
  assign n8471 = n8470 ^ n6419 ;
  assign n8472 = n8471 ^ n6222 ;
  assign n8482 = n8481 ^ n8472 ;
  assign n8484 = n8482 ^ x437 ;
  assign n8483 = n8482 ^ n8461 ;
  assign n8485 = n8484 ^ n8483 ;
  assign n8486 = n8466 & ~n8485 ;
  assign n8487 = n8486 ^ n8484 ;
  assign n8500 = n7922 ^ n7921 ;
  assign n8496 = n7694 ^ n7686 ;
  assign n8495 = n8478 ^ n7694 ;
  assign n8497 = n8496 ^ n8495 ;
  assign n8498 = ~n8477 & n8497 ;
  assign n8499 = n8498 ^ n8496 ;
  assign n8501 = n8500 ^ n8499 ;
  assign n8502 = ~n7502 & ~n8501 ;
  assign n8503 = n8502 ^ n7145 ;
  assign n8490 = n8481 ^ n8471 ;
  assign n8491 = n8481 ^ n6222 ;
  assign n8492 = ~n8490 & n8491 ;
  assign n8493 = n8492 ^ n6222 ;
  assign n8494 = n8493 ^ n6434 ;
  assign n8504 = n8503 ^ n8494 ;
  assign n8506 = n8504 ^ x436 ;
  assign n8505 = n8504 ^ n8482 ;
  assign n8507 = n8506 ^ n8505 ;
  assign n8508 = n8487 & ~n8507 ;
  assign n8509 = n8508 ^ n8506 ;
  assign n8510 = n8509 ^ x435 ;
  assign n8025 = n8024 ^ x421 ;
  assign n8026 = n7981 ^ x423 ;
  assign n8027 = n7982 ^ x422 ;
  assign n8028 = n8027 ^ n7980 ;
  assign n8029 = n8026 & n8028 ;
  assign n8030 = ~n8025 & ~n8029 ;
  assign n8072 = n8071 ^ x420 ;
  assign n8073 = n8030 & n8072 ;
  assign n8116 = n8115 ^ x419 ;
  assign n8117 = ~n8073 & ~n8116 ;
  assign n8159 = n8158 ^ x418 ;
  assign n8160 = ~n8117 & n8159 ;
  assign n8201 = n8200 ^ x417 ;
  assign n8202 = n8160 & n8201 ;
  assign n8224 = n8223 ^ x416 ;
  assign n8225 = ~n8202 & ~n8224 ;
  assign n8239 = n8238 ^ x431 ;
  assign n8243 = n8242 ^ n8239 ;
  assign n8244 = n8225 & ~n8243 ;
  assign n8267 = n8266 ^ x430 ;
  assign n8268 = ~n8244 & n8267 ;
  assign n8289 = n8288 ^ x429 ;
  assign n8290 = n8268 & n8289 ;
  assign n8312 = n8311 ^ x428 ;
  assign n8313 = n8290 & ~n8312 ;
  assign n8333 = n8332 ^ x427 ;
  assign n8334 = ~n8313 & n8333 ;
  assign n8355 = n8354 ^ x426 ;
  assign n8356 = n8334 & n8355 ;
  assign n8378 = n8377 ^ x425 ;
  assign n8379 = n8356 & ~n8378 ;
  assign n8399 = n8398 ^ x424 ;
  assign n8400 = ~n8379 & n8399 ;
  assign n8422 = n8421 ^ x439 ;
  assign n8423 = n8400 & ~n8422 ;
  assign n8444 = n8443 ^ x438 ;
  assign n8445 = n8423 & n8444 ;
  assign n8467 = n8466 ^ x437 ;
  assign n8468 = n8445 & ~n8467 ;
  assign n8488 = n8487 ^ x436 ;
  assign n8489 = ~n8468 & n8488 ;
  assign n8511 = n8510 ^ n8489 ;
  assign n9090 = n8520 ^ n8511 ;
  assign n8534 = n7924 ^ n7923 ;
  assign n8530 = n7703 ^ n7694 ;
  assign n8529 = n8500 ^ n7703 ;
  assign n8531 = n8530 ^ n8529 ;
  assign n8532 = n8499 & n8531 ;
  assign n8533 = n8532 ^ n8530 ;
  assign n8535 = n8534 ^ n8533 ;
  assign n8536 = n7527 & n8535 ;
  assign n8537 = n8536 ^ n7156 ;
  assign n8524 = n8503 ^ n8493 ;
  assign n8525 = n8503 ^ n6434 ;
  assign n8526 = n8524 & n8525 ;
  assign n8527 = n8526 ^ n6434 ;
  assign n8528 = n8527 ^ n6442 ;
  assign n8538 = n8537 ^ n8528 ;
  assign n8540 = n8538 ^ x435 ;
  assign n8539 = n8538 ^ n8504 ;
  assign n8541 = n8540 ^ n8539 ;
  assign n8542 = n8509 & ~n8541 ;
  assign n8543 = n8542 ^ n8540 ;
  assign n8544 = n8543 ^ x434 ;
  assign n8523 = n8489 & n8510 ;
  assign n8545 = n8544 ^ n8523 ;
  assign n8521 = ~n8511 & n8520 ;
  assign n8522 = n8521 ^ n7977 ;
  assign n8546 = n8545 ^ n8522 ;
  assign n8547 = ~n8012 & n8546 ;
  assign n8548 = n8547 ^ n7595 ;
  assign n8512 = n8511 ^ n7974 ;
  assign n8513 = n7946 & n8512 ;
  assign n8514 = n8513 ^ n7974 ;
  assign n8518 = ~n7395 & n8514 ;
  assign n8519 = n8518 ^ n6885 ;
  assign n8549 = n8548 ^ n8519 ;
  assign n8515 = n8514 ^ n7395 ;
  assign n8516 = x455 & ~n8515 ;
  assign n8551 = n8549 ^ n8516 ;
  assign n8568 = n7711 ^ n7175 ;
  assign n8574 = n7926 ^ n7925 ;
  assign n8570 = n7711 ^ n7703 ;
  assign n8569 = n8534 ^ n7711 ;
  assign n8571 = n8570 ^ n8569 ;
  assign n8572 = ~n8533 & ~n8571 ;
  assign n8573 = n8572 ^ n8570 ;
  assign n8575 = n8574 ^ n8573 ;
  assign n8576 = ~n8568 & ~n8575 ;
  assign n8577 = n8576 ^ n7175 ;
  assign n8563 = n8537 ^ n8527 ;
  assign n8564 = n8537 ^ n6442 ;
  assign n8565 = ~n8563 & n8564 ;
  assign n8566 = n8565 ^ n6442 ;
  assign n8567 = n8566 ^ n6450 ;
  assign n8578 = n8577 ^ n8567 ;
  assign n8580 = n8578 ^ x434 ;
  assign n8579 = n8578 ^ n8538 ;
  assign n8581 = n8580 ^ n8579 ;
  assign n8582 = ~n8543 & n8581 ;
  assign n8583 = n8582 ^ n8580 ;
  assign n8584 = n8583 ^ x433 ;
  assign n8562 = ~n8523 & n8544 ;
  assign n8585 = n8584 ^ n8562 ;
  assign n8557 = n8545 ^ n8521 ;
  assign n8558 = n8545 ^ n7977 ;
  assign n8559 = n8557 & n8558 ;
  assign n8560 = n8559 ^ n7977 ;
  assign n8561 = n8560 ^ n8016 ;
  assign n8586 = n8585 ^ n8561 ;
  assign n8587 = n8035 & n8586 ;
  assign n8588 = n8587 ^ n7592 ;
  assign n8552 = n8548 ^ n8518 ;
  assign n8553 = n8548 ^ n6885 ;
  assign n8554 = ~n8552 & ~n8553 ;
  assign n8555 = n8554 ^ n6885 ;
  assign n8556 = n8555 ^ n6892 ;
  assign n8589 = n8588 ^ n8556 ;
  assign n8590 = n8589 ^ x454 ;
  assign n8591 = n8590 ^ n8549 ;
  assign n8592 = n8591 ^ n8589 ;
  assign n8593 = n8551 & ~n8592 ;
  assign n8594 = n8593 ^ n8590 ;
  assign n8626 = n8585 ^ n8560 ;
  assign n8627 = n8585 ^ n8016 ;
  assign n8628 = ~n8626 & ~n8627 ;
  assign n8629 = n8628 ^ n8016 ;
  assign n8630 = n8629 ^ n8063 ;
  assign n8608 = n7539 ^ n6869 ;
  assign n8614 = n7928 ^ n7927 ;
  assign n8610 = n7711 ^ n7539 ;
  assign n8609 = n8574 ^ n7539 ;
  assign n8611 = n8610 ^ n8609 ;
  assign n8612 = n8573 & ~n8611 ;
  assign n8613 = n8612 ^ n8610 ;
  assign n8615 = n8614 ^ n8613 ;
  assign n8616 = n8608 & ~n8615 ;
  assign n8617 = n8616 ^ n6869 ;
  assign n8603 = n8577 ^ n8566 ;
  assign n8604 = n8577 ^ n6450 ;
  assign n8605 = n8603 & ~n8604 ;
  assign n8606 = n8605 ^ n6450 ;
  assign n8607 = n8606 ^ n6458 ;
  assign n8618 = n8617 ^ n8607 ;
  assign n8620 = n8618 ^ x433 ;
  assign n8619 = n8618 ^ n8578 ;
  assign n8621 = n8620 ^ n8619 ;
  assign n8622 = n8583 & ~n8621 ;
  assign n8623 = n8622 ^ n8620 ;
  assign n8624 = n8623 ^ x432 ;
  assign n8602 = n8562 & ~n8584 ;
  assign n8625 = n8624 ^ n8602 ;
  assign n8631 = n8630 ^ n8625 ;
  assign n8632 = n8103 & ~n8631 ;
  assign n8633 = n8632 ^ n7589 ;
  assign n8597 = n8588 ^ n8555 ;
  assign n8598 = n8588 ^ n6892 ;
  assign n8599 = n8597 & n8598 ;
  assign n8600 = n8599 ^ n6892 ;
  assign n8601 = n8600 ^ n6900 ;
  assign n8634 = n8633 ^ n8601 ;
  assign n8636 = n8634 ^ x453 ;
  assign n8635 = n8634 ^ n8589 ;
  assign n8637 = n8636 ^ n8635 ;
  assign n8638 = n8594 & ~n8637 ;
  assign n8639 = n8638 ^ n8636 ;
  assign n8653 = n8617 ^ n8606 ;
  assign n8659 = n7930 ^ n7929 ;
  assign n8655 = n7724 ^ n7539 ;
  assign n8654 = n8614 ^ n7724 ;
  assign n8656 = n8655 ^ n8654 ;
  assign n8657 = n8613 & ~n8656 ;
  assign n8658 = n8657 ^ n8655 ;
  assign n8660 = n8659 ^ n8658 ;
  assign n8661 = ~n7875 & ~n8660 ;
  assign n8662 = n8661 ^ n7206 ;
  assign n8663 = n8662 ^ n6458 ;
  assign n8664 = n8663 ^ n8662 ;
  assign n8665 = n8664 ^ n8606 ;
  assign n8666 = ~n8653 & ~n8665 ;
  assign n8667 = n8666 ^ n8663 ;
  assign n8668 = n8667 ^ n6463 ;
  assign n8670 = n8668 ^ x432 ;
  assign n8669 = n8668 ^ n8618 ;
  assign n8671 = n8670 ^ n8669 ;
  assign n8672 = n8623 & ~n8671 ;
  assign n8673 = n8672 ^ n8670 ;
  assign n8674 = n8673 ^ x447 ;
  assign n8652 = ~n8602 & n8624 ;
  assign n8675 = n8674 ^ n8652 ;
  assign n8647 = n8625 ^ n8063 ;
  assign n8648 = n8629 ^ n8625 ;
  assign n8649 = ~n8647 & ~n8648 ;
  assign n8650 = n8649 ^ n8063 ;
  assign n8651 = n8650 ^ n8107 ;
  assign n8676 = n8675 ^ n8651 ;
  assign n8677 = n8122 & ~n8676 ;
  assign n8678 = n8677 ^ n7585 ;
  assign n8642 = n8633 ^ n8600 ;
  assign n8643 = n8633 ^ n6900 ;
  assign n8644 = n8642 & n8643 ;
  assign n8645 = n8644 ^ n6900 ;
  assign n8646 = n8645 ^ n6907 ;
  assign n8679 = n8678 ^ n8646 ;
  assign n8681 = n8679 ^ x452 ;
  assign n8680 = n8679 ^ n8634 ;
  assign n8682 = n8681 ^ n8680 ;
  assign n8683 = ~n8639 & n8682 ;
  assign n8684 = n8683 ^ n8681 ;
  assign n8714 = n8675 ^ n8650 ;
  assign n8715 = n8675 ^ n8107 ;
  assign n8716 = ~n8714 & n8715 ;
  assign n8717 = n8716 ^ n8107 ;
  assign n8718 = n8717 ^ n8150 ;
  assign n8697 = n7883 ^ n7876 ;
  assign n8699 = n8659 ^ n7724 ;
  assign n8700 = ~n8658 & ~n8699 ;
  assign n8701 = n8700 ^ n7724 ;
  assign n8698 = n7932 ^ n7931 ;
  assign n8702 = n8701 ^ n8698 ;
  assign n8703 = n8702 ^ n7883 ;
  assign n8704 = ~n8697 & ~n8703 ;
  assign n8705 = n8704 ^ n7876 ;
  assign n8693 = n8662 ^ n6463 ;
  assign n8694 = n8667 & n8693 ;
  assign n8695 = n8694 ^ n6463 ;
  assign n8696 = n8695 ^ n7240 ;
  assign n8706 = n8705 ^ n8696 ;
  assign n8708 = n8706 ^ x447 ;
  assign n8707 = n8706 ^ n8668 ;
  assign n8709 = n8708 ^ n8707 ;
  assign n8710 = n8673 & ~n8709 ;
  assign n8711 = n8710 ^ n8708 ;
  assign n8712 = n8711 ^ x446 ;
  assign n8692 = n8652 & n8674 ;
  assign n8713 = n8712 ^ n8692 ;
  assign n8719 = n8718 ^ n8713 ;
  assign n8720 = ~n8165 & ~n8719 ;
  assign n8721 = n8720 ^ n7582 ;
  assign n8687 = n8678 ^ n8645 ;
  assign n8688 = n8678 ^ n6907 ;
  assign n8689 = ~n8687 & n8688 ;
  assign n8690 = n8689 ^ n6907 ;
  assign n8691 = n8690 ^ n6915 ;
  assign n8722 = n8721 ^ n8691 ;
  assign n8724 = n8722 ^ x451 ;
  assign n8723 = n8722 ^ n8679 ;
  assign n8725 = n8724 ^ n8723 ;
  assign n8726 = n8684 & ~n8725 ;
  assign n8727 = n8726 ^ n8724 ;
  assign n8745 = n7962 ^ n7246 ;
  assign n8751 = n7934 ^ n7933 ;
  assign n8747 = n7962 ^ n7883 ;
  assign n8746 = n8701 ^ n7962 ;
  assign n8748 = n8747 ^ n8746 ;
  assign n8749 = n8702 & ~n8748 ;
  assign n8750 = n8749 ^ n8747 ;
  assign n8752 = n8751 ^ n8750 ;
  assign n8753 = ~n8745 & n8752 ;
  assign n8754 = n8753 ^ n7246 ;
  assign n8740 = n8705 ^ n8695 ;
  assign n8741 = n8705 ^ n7240 ;
  assign n8742 = n8740 & ~n8741 ;
  assign n8743 = n8742 ^ n7240 ;
  assign n8744 = n8743 ^ n6298 ;
  assign n8755 = n8754 ^ n8744 ;
  assign n8757 = n8755 ^ x446 ;
  assign n8756 = n8755 ^ n8706 ;
  assign n8758 = n8757 ^ n8756 ;
  assign n8759 = n8711 & ~n8758 ;
  assign n8760 = n8759 ^ n8757 ;
  assign n8761 = n8760 ^ x445 ;
  assign n8739 = ~n8692 & ~n8712 ;
  assign n8762 = n8761 ^ n8739 ;
  assign n8763 = n8762 ^ n8192 ;
  assign n8735 = n8713 ^ n8150 ;
  assign n8736 = n8717 ^ n8713 ;
  assign n8737 = n8735 & n8736 ;
  assign n8738 = n8737 ^ n8150 ;
  assign n8764 = n8763 ^ n8738 ;
  assign n8765 = ~n8208 & n8764 ;
  assign n8766 = n8765 ^ n7578 ;
  assign n8730 = n8721 ^ n8690 ;
  assign n8731 = n8721 ^ n6915 ;
  assign n8732 = ~n8730 & ~n8731 ;
  assign n8733 = n8732 ^ n6915 ;
  assign n8734 = n8733 ^ n6922 ;
  assign n8767 = n8766 ^ n8734 ;
  assign n8769 = n8767 ^ x450 ;
  assign n8768 = n8767 ^ n8722 ;
  assign n8770 = n8769 ^ n8768 ;
  assign n8771 = ~n8727 & n8770 ;
  assign n8772 = n8771 ^ n8769 ;
  assign n8780 = n8215 ^ n7575 ;
  assign n8805 = n8762 ^ n8738 ;
  assign n8806 = n8763 & ~n8805 ;
  assign n8807 = n8806 ^ n8192 ;
  assign n8808 = n8807 ^ n8215 ;
  assign n8787 = n8000 ^ n7267 ;
  assign n8793 = n7936 ^ n7935 ;
  assign n8789 = n8000 ^ n7962 ;
  assign n8788 = n8751 ^ n8000 ;
  assign n8790 = n8789 ^ n8788 ;
  assign n8791 = ~n8750 & n8790 ;
  assign n8792 = n8791 ^ n8789 ;
  assign n8794 = n8793 ^ n8792 ;
  assign n8795 = n8787 & ~n8794 ;
  assign n8796 = n8795 ^ n7267 ;
  assign n8782 = n8754 ^ n8743 ;
  assign n8783 = n8754 ^ n6298 ;
  assign n8784 = ~n8782 & ~n8783 ;
  assign n8785 = n8784 ^ n6298 ;
  assign n8786 = n8785 ^ n7260 ;
  assign n8797 = n8796 ^ n8786 ;
  assign n8799 = n8797 ^ x445 ;
  assign n8798 = n8797 ^ n8755 ;
  assign n8800 = n8799 ^ n8798 ;
  assign n8801 = n8760 & ~n8800 ;
  assign n8802 = n8801 ^ n8799 ;
  assign n8803 = n8802 ^ x444 ;
  assign n8781 = ~n8739 & n8761 ;
  assign n8804 = n8803 ^ n8781 ;
  assign n8809 = n8808 ^ n8804 ;
  assign n8810 = ~n8780 & n8809 ;
  assign n8811 = n8810 ^ n7575 ;
  assign n8775 = n8766 ^ n8733 ;
  assign n8776 = n8766 ^ n6922 ;
  assign n8777 = n8775 & n8776 ;
  assign n8778 = n8777 ^ n6922 ;
  assign n8779 = n8778 ^ n6930 ;
  assign n8812 = n8811 ^ n8779 ;
  assign n8814 = n8812 ^ x449 ;
  assign n8813 = n8812 ^ n8767 ;
  assign n8815 = n8814 ^ n8813 ;
  assign n8816 = ~n8772 & n8815 ;
  assign n8817 = n8816 ^ n8814 ;
  assign n8835 = n8051 ^ n7291 ;
  assign n8841 = n7938 ^ n7937 ;
  assign n8837 = n8051 ^ n8000 ;
  assign n8836 = n8793 ^ n8051 ;
  assign n8838 = n8837 ^ n8836 ;
  assign n8839 = n8792 & n8838 ;
  assign n8840 = n8839 ^ n8837 ;
  assign n8842 = n8841 ^ n8840 ;
  assign n8843 = n8835 & ~n8842 ;
  assign n8844 = n8843 ^ n7291 ;
  assign n8830 = n8796 ^ n8785 ;
  assign n8831 = n8796 ^ n7260 ;
  assign n8832 = ~n8830 & ~n8831 ;
  assign n8833 = n8832 ^ n7260 ;
  assign n8834 = n8833 ^ n6494 ;
  assign n8845 = n8844 ^ n8834 ;
  assign n8847 = n8845 ^ x444 ;
  assign n8846 = n8845 ^ n8797 ;
  assign n8848 = n8847 ^ n8846 ;
  assign n8849 = ~n8802 & n8848 ;
  assign n8850 = n8849 ^ n8847 ;
  assign n8851 = n8850 ^ x443 ;
  assign n8829 = n8781 & ~n8803 ;
  assign n8852 = n8851 ^ n8829 ;
  assign n8825 = n8807 ^ n8804 ;
  assign n8826 = n8808 & ~n8825 ;
  assign n8827 = n8826 ^ n8215 ;
  assign n8828 = n8827 ^ n8235 ;
  assign n8853 = n8852 ^ n8828 ;
  assign n8854 = ~n8251 & ~n8853 ;
  assign n8855 = n8854 ^ n7572 ;
  assign n8820 = n8811 ^ n8778 ;
  assign n8821 = n8811 ^ n6930 ;
  assign n8822 = ~n8820 & n8821 ;
  assign n8823 = n8822 ^ n6930 ;
  assign n8824 = n8823 ^ n6937 ;
  assign n8856 = n8855 ^ n8824 ;
  assign n8858 = n8856 ^ x448 ;
  assign n8857 = n8856 ^ n8812 ;
  assign n8859 = n8858 ^ n8857 ;
  assign n8860 = n8817 & ~n8859 ;
  assign n8861 = n8860 ^ n8858 ;
  assign n8869 = n8258 ^ n7568 ;
  assign n8894 = n8852 ^ n8827 ;
  assign n8895 = n8852 ^ n8235 ;
  assign n8896 = ~n8894 & ~n8895 ;
  assign n8897 = n8896 ^ n8235 ;
  assign n8898 = n8897 ^ n8258 ;
  assign n8876 = n8090 ^ n7312 ;
  assign n8882 = n7940 ^ n7939 ;
  assign n8878 = n8090 ^ n8051 ;
  assign n8877 = n8841 ^ n8090 ;
  assign n8879 = n8878 ^ n8877 ;
  assign n8880 = ~n8840 & n8879 ;
  assign n8881 = n8880 ^ n8878 ;
  assign n8883 = n8882 ^ n8881 ;
  assign n8884 = ~n8876 & ~n8883 ;
  assign n8885 = n8884 ^ n7312 ;
  assign n8871 = n8844 ^ n8833 ;
  assign n8872 = n8844 ^ n6494 ;
  assign n8873 = ~n8871 & n8872 ;
  assign n8874 = n8873 ^ n6494 ;
  assign n8875 = n8874 ^ n6502 ;
  assign n8886 = n8885 ^ n8875 ;
  assign n8888 = n8886 ^ x443 ;
  assign n8887 = n8886 ^ n8845 ;
  assign n8889 = n8888 ^ n8887 ;
  assign n8890 = ~n8850 & n8889 ;
  assign n8891 = n8890 ^ n8888 ;
  assign n8892 = n8891 ^ x442 ;
  assign n8870 = n8829 & ~n8851 ;
  assign n8893 = n8892 ^ n8870 ;
  assign n8899 = n8898 ^ n8893 ;
  assign n8900 = ~n8869 & ~n8899 ;
  assign n8901 = n8900 ^ n7568 ;
  assign n8864 = n8855 ^ n8823 ;
  assign n8865 = n8855 ^ n6937 ;
  assign n8866 = n8864 & n8865 ;
  assign n8867 = n8866 ^ n6937 ;
  assign n8868 = n8867 ^ n6945 ;
  assign n8902 = n8901 ^ n8868 ;
  assign n8904 = n8902 ^ x463 ;
  assign n8903 = n8902 ^ n8856 ;
  assign n8905 = n8904 ^ n8903 ;
  assign n8906 = n8861 & ~n8905 ;
  assign n8907 = n8906 ^ n8904 ;
  assign n8915 = n8280 ^ n7564 ;
  assign n8927 = n8139 ^ n7490 ;
  assign n8933 = n7942 ^ n7941 ;
  assign n8929 = n8139 ^ n8090 ;
  assign n8928 = n8882 ^ n8139 ;
  assign n8930 = n8929 ^ n8928 ;
  assign n8931 = n8881 & ~n8930 ;
  assign n8932 = n8931 ^ n8929 ;
  assign n8934 = n8933 ^ n8932 ;
  assign n8935 = ~n8927 & ~n8934 ;
  assign n8936 = n8935 ^ n7490 ;
  assign n8922 = n8885 ^ n8874 ;
  assign n8923 = n8885 ^ n6502 ;
  assign n8924 = n8922 & n8923 ;
  assign n8925 = n8924 ^ n6502 ;
  assign n8926 = n8925 ^ n6510 ;
  assign n8937 = n8936 ^ n8926 ;
  assign n8939 = n8937 ^ x442 ;
  assign n8938 = n8937 ^ n8886 ;
  assign n8940 = n8939 ^ n8938 ;
  assign n8941 = ~n8891 & n8940 ;
  assign n8942 = n8941 ^ n8939 ;
  assign n8943 = n8942 ^ x441 ;
  assign n8921 = n8870 & ~n8892 ;
  assign n8944 = n8943 ^ n8921 ;
  assign n8916 = n8893 ^ n8258 ;
  assign n8917 = n8897 ^ n8893 ;
  assign n8918 = n8916 & n8917 ;
  assign n8919 = n8918 ^ n8258 ;
  assign n8920 = n8919 ^ n8280 ;
  assign n8945 = n8944 ^ n8920 ;
  assign n8946 = n8915 & n8945 ;
  assign n8947 = n8946 ^ n7564 ;
  assign n8910 = n8901 ^ n8867 ;
  assign n8911 = n8901 ^ n6945 ;
  assign n8912 = n8910 & n8911 ;
  assign n8913 = n8912 ^ n6945 ;
  assign n8914 = n8913 ^ n6952 ;
  assign n8948 = n8947 ^ n8914 ;
  assign n8950 = n8948 ^ x462 ;
  assign n8949 = n8948 ^ n8902 ;
  assign n8951 = n8950 ^ n8949 ;
  assign n8952 = ~n8907 & n8951 ;
  assign n8953 = n8952 ^ n8950 ;
  assign n8983 = n8944 ^ n8919 ;
  assign n8984 = n8944 ^ n8280 ;
  assign n8985 = ~n8983 & n8984 ;
  assign n8986 = n8985 ^ n8280 ;
  assign n8987 = n8986 ^ n8298 ;
  assign n8973 = n8187 ^ n7515 ;
  assign n8977 = n8933 ^ n8139 ;
  assign n8978 = ~n8932 & ~n8977 ;
  assign n8974 = n7944 ^ n7943 ;
  assign n8975 = n8974 ^ n8187 ;
  assign n8976 = n8975 ^ n8933 ;
  assign n8979 = n8978 ^ n8976 ;
  assign n8980 = ~n8973 & ~n8979 ;
  assign n8970 = n6510 ^ x440 ;
  assign n8971 = n8970 ^ n8181 ;
  assign n8967 = n8936 ^ n8925 ;
  assign n8968 = n8936 ^ n6510 ;
  assign n8969 = ~n8967 & ~n8968 ;
  assign n8972 = n8971 ^ n8969 ;
  assign n8981 = n8980 ^ n8972 ;
  assign n8962 = n8937 ^ n8921 ;
  assign n8965 = ~n8942 & n8962 ;
  assign n8961 = n8942 ^ n8937 ;
  assign n8963 = n8962 ^ n8961 ;
  assign n8964 = x441 & n8963 ;
  assign n8966 = n8965 ^ n8964 ;
  assign n8982 = n8981 ^ n8966 ;
  assign n8988 = n8987 ^ n8982 ;
  assign n8989 = ~n8297 & n8988 ;
  assign n8990 = n8989 ^ n7561 ;
  assign n8956 = n8947 ^ n8913 ;
  assign n8957 = n8947 ^ n6952 ;
  assign n8958 = n8956 & ~n8957 ;
  assign n8959 = n8958 ^ n6952 ;
  assign n8960 = n8959 ^ n6877 ;
  assign n8991 = n8990 ^ n8960 ;
  assign n8993 = n8991 ^ x461 ;
  assign n8992 = n8991 ^ n8948 ;
  assign n8994 = n8993 ^ n8992 ;
  assign n8995 = ~n8953 & n8994 ;
  assign n8996 = n8995 ^ n8993 ;
  assign n9008 = n8990 ^ n8959 ;
  assign n9009 = n8990 ^ n6877 ;
  assign n9010 = n9008 & ~n9009 ;
  assign n9011 = n9010 ^ n6877 ;
  assign n9012 = n9011 ^ n6872 ;
  assign n8999 = n8324 ^ n7557 ;
  assign n9004 = n8324 ^ n8026 ;
  assign n9000 = n8982 ^ n8298 ;
  assign n9001 = n8986 ^ n8982 ;
  assign n9002 = n9000 & n9001 ;
  assign n9003 = n9002 ^ n8298 ;
  assign n9005 = n9004 ^ n9003 ;
  assign n9006 = ~n8999 & n9005 ;
  assign n9007 = n9006 ^ n7557 ;
  assign n9013 = n9012 ^ n9007 ;
  assign n9015 = n9013 ^ x460 ;
  assign n9014 = n9013 ^ n8991 ;
  assign n9016 = n9015 ^ n9014 ;
  assign n9017 = ~n8996 & n9016 ;
  assign n9018 = n9017 ^ n9015 ;
  assign n9032 = n9011 ^ n9007 ;
  assign n9033 = n9007 ^ n6872 ;
  assign n9034 = n9032 & n9033 ;
  assign n9035 = n9034 ^ n6872 ;
  assign n9036 = n9035 ^ n6967 ;
  assign n9021 = n8346 ^ n7554 ;
  assign n9028 = n8028 ^ n8026 ;
  assign n9022 = n9003 ^ n8026 ;
  assign n9023 = n8346 ^ n8324 ;
  assign n9024 = n9023 ^ n8346 ;
  assign n9025 = n9024 ^ n9003 ;
  assign n9026 = n9022 & n9025 ;
  assign n9027 = n9026 ^ n9023 ;
  assign n9029 = n9028 ^ n9027 ;
  assign n9030 = ~n9021 & n9029 ;
  assign n9031 = n9030 ^ n7554 ;
  assign n9037 = n9036 ^ n9031 ;
  assign n9039 = n9037 ^ x459 ;
  assign n9038 = n9037 ^ n9013 ;
  assign n9040 = n9039 ^ n9038 ;
  assign n9041 = n9018 & ~n9040 ;
  assign n9042 = n9041 ^ n9039 ;
  assign n9050 = n8364 ^ n7550 ;
  assign n9056 = n8029 ^ n8025 ;
  assign n9052 = n8364 ^ n8346 ;
  assign n9051 = n9028 ^ n8364 ;
  assign n9053 = n9052 ^ n9051 ;
  assign n9054 = ~n9027 & ~n9053 ;
  assign n9055 = n9054 ^ n9052 ;
  assign n9057 = n9056 ^ n9055 ;
  assign n9058 = ~n9050 & ~n9057 ;
  assign n9059 = n9058 ^ n7550 ;
  assign n9045 = n9031 ^ n6967 ;
  assign n9046 = n9035 ^ n9031 ;
  assign n9047 = ~n9045 & n9046 ;
  assign n9048 = n9047 ^ n6967 ;
  assign n9049 = n9048 ^ n6977 ;
  assign n9060 = n9059 ^ n9049 ;
  assign n9062 = n9060 ^ x458 ;
  assign n9061 = n9060 ^ n9037 ;
  assign n9063 = n9062 ^ n9061 ;
  assign n9064 = n9042 & ~n9063 ;
  assign n9065 = n9064 ^ n9062 ;
  assign n9077 = n9059 ^ n9048 ;
  assign n9078 = n9059 ^ n6977 ;
  assign n9079 = ~n9077 & ~n9078 ;
  assign n9080 = n9079 ^ n6977 ;
  assign n9081 = n9080 ^ n7070 ;
  assign n9068 = n8390 ^ n7547 ;
  assign n9070 = n9056 ^ n8364 ;
  assign n9071 = ~n9055 & ~n9070 ;
  assign n9072 = n9071 ^ n8364 ;
  assign n9069 = n8072 ^ n8030 ;
  assign n9073 = n9072 ^ n9069 ;
  assign n9074 = n9073 ^ n8390 ;
  assign n9075 = n9068 & ~n9074 ;
  assign n9076 = n9075 ^ n7547 ;
  assign n9082 = n9081 ^ n9076 ;
  assign n9084 = n9082 ^ x457 ;
  assign n9083 = n9082 ^ n9060 ;
  assign n9085 = n9084 ^ n9083 ;
  assign n9086 = n9065 & ~n9085 ;
  assign n9087 = n9086 ^ n9084 ;
  assign n9088 = n9087 ^ x456 ;
  assign n8517 = n8516 ^ x454 ;
  assign n8550 = n8549 ^ n8517 ;
  assign n8595 = n8594 ^ x453 ;
  assign n8596 = n8550 & n8595 ;
  assign n8640 = n8639 ^ x452 ;
  assign n8641 = n8596 & ~n8640 ;
  assign n8685 = n8684 ^ x451 ;
  assign n8686 = ~n8641 & ~n8685 ;
  assign n8728 = n8727 ^ x450 ;
  assign n8729 = n8686 & n8728 ;
  assign n8773 = n8772 ^ x449 ;
  assign n8774 = n8729 & n8773 ;
  assign n8818 = n8817 ^ x448 ;
  assign n8819 = ~n8774 & n8818 ;
  assign n8862 = n8861 ^ x463 ;
  assign n8863 = n8819 & n8862 ;
  assign n8908 = n8907 ^ x462 ;
  assign n8909 = n8863 & ~n8908 ;
  assign n8954 = n8953 ^ x461 ;
  assign n8955 = ~n8909 & n8954 ;
  assign n8997 = n8996 ^ x460 ;
  assign n8998 = n8955 & n8997 ;
  assign n9019 = n9018 ^ x459 ;
  assign n9020 = n8998 & ~n9019 ;
  assign n9043 = n9042 ^ x458 ;
  assign n9044 = n9020 & ~n9043 ;
  assign n9066 = n9065 ^ x457 ;
  assign n9067 = ~n9044 & n9066 ;
  assign n9089 = n9088 ^ n9067 ;
  assign n9091 = n9090 ^ n9089 ;
  assign n9555 = n8378 ^ n8356 ;
  assign n9106 = n8408 ^ n8390 ;
  assign n9105 = n9072 ^ n8408 ;
  assign n9107 = n9106 ^ n9105 ;
  assign n9108 = n9073 & ~n9107 ;
  assign n9109 = n9108 ^ n9106 ;
  assign n9110 = n8116 ^ n8073 ;
  assign n9147 = n9110 ^ n8408 ;
  assign n9148 = ~n9109 & n9147 ;
  assign n9149 = n9148 ^ n8408 ;
  assign n9193 = n9149 ^ n8453 ;
  assign n9146 = n8159 ^ n8117 ;
  assign n9150 = n9149 ^ n9146 ;
  assign n9190 = n8434 ^ n7542 ;
  assign n9191 = n9190 ^ n9149 ;
  assign n9192 = n9150 & n9191 ;
  assign n9194 = n9193 ^ n9192 ;
  assign n9240 = n8479 ^ n8453 ;
  assign n9195 = n8201 ^ n8160 ;
  assign n9239 = n9195 ^ n8479 ;
  assign n9241 = n9240 ^ n9239 ;
  assign n9242 = n9194 & ~n9241 ;
  assign n9243 = n9242 ^ n9240 ;
  assign n9285 = n8501 ^ n8479 ;
  assign n9244 = n8224 ^ n8202 ;
  assign n9284 = n9244 ^ n8501 ;
  assign n9286 = n9285 ^ n9284 ;
  assign n9287 = ~n9243 & ~n9286 ;
  assign n9288 = n9287 ^ n9285 ;
  assign n9330 = n8535 ^ n8501 ;
  assign n9289 = n8243 ^ n8225 ;
  assign n9329 = n9289 ^ n8535 ;
  assign n9331 = n9330 ^ n9329 ;
  assign n9332 = ~n9288 & ~n9331 ;
  assign n9333 = n9332 ^ n9330 ;
  assign n9375 = n8575 ^ n8535 ;
  assign n9334 = n8267 ^ n8244 ;
  assign n9374 = n9334 ^ n8575 ;
  assign n9376 = n9375 ^ n9374 ;
  assign n9377 = ~n9333 & ~n9376 ;
  assign n9378 = n9377 ^ n9375 ;
  assign n9420 = n8615 ^ n8575 ;
  assign n9379 = n8289 ^ n8268 ;
  assign n9419 = n9379 ^ n8615 ;
  assign n9421 = n9420 ^ n9419 ;
  assign n9422 = ~n9378 & ~n9421 ;
  assign n9423 = n9422 ^ n9420 ;
  assign n9464 = n8660 ^ n8615 ;
  assign n9424 = n8312 ^ n8290 ;
  assign n9463 = n9424 ^ n8660 ;
  assign n9465 = n9464 ^ n9463 ;
  assign n9466 = n9423 & n9465 ;
  assign n9467 = n9466 ^ n9464 ;
  assign n9468 = n8333 ^ n8313 ;
  assign n9503 = n9468 ^ n8660 ;
  assign n9504 = n9467 & ~n9503 ;
  assign n9505 = n9504 ^ n8660 ;
  assign n9502 = n8355 ^ n8334 ;
  assign n9506 = n9505 ^ n9502 ;
  assign n9551 = n8752 ^ n8703 ;
  assign n9550 = n9505 ^ n8752 ;
  assign n9552 = n9551 ^ n9550 ;
  assign n9553 = ~n9506 & n9552 ;
  assign n9554 = n9553 ^ n9551 ;
  assign n9556 = n9555 ^ n9554 ;
  assign n9104 = n9080 ^ n9076 ;
  assign n9111 = n9110 ^ n9109 ;
  assign n9112 = n8408 ^ n7660 ;
  assign n9113 = n9111 & ~n9112 ;
  assign n9114 = n9113 ^ n7660 ;
  assign n9115 = n9114 ^ n7070 ;
  assign n9116 = n9115 ^ n9114 ;
  assign n9117 = n9116 ^ n9080 ;
  assign n9118 = n9104 & ~n9117 ;
  assign n9119 = n9118 ^ n9115 ;
  assign n9120 = n9119 ^ n7081 ;
  assign n9122 = n9120 ^ x456 ;
  assign n9121 = n9120 ^ n9082 ;
  assign n9123 = n9122 ^ n9121 ;
  assign n9124 = n9087 & ~n9123 ;
  assign n9125 = n9124 ^ n9122 ;
  assign n9126 = n9125 ^ x471 ;
  assign n9103 = ~n9067 & ~n9088 ;
  assign n9127 = n9126 ^ n9103 ;
  assign n9101 = n9089 & ~n9090 ;
  assign n9102 = n9101 ^ n8546 ;
  assign n9128 = n9127 ^ n9102 ;
  assign n9129 = ~n8557 & n9128 ;
  assign n9130 = n9129 ^ n7977 ;
  assign n9092 = n9089 ^ n8520 ;
  assign n9093 = ~n8511 & ~n9092 ;
  assign n9094 = n9093 ^ n8520 ;
  assign n9099 = n7974 & n9094 ;
  assign n9100 = n9099 ^ n7595 ;
  assign n9131 = n9130 ^ n9100 ;
  assign n9095 = n9094 ^ n7974 ;
  assign n9097 = x487 & n9095 ;
  assign n9134 = n9131 ^ n9097 ;
  assign n9154 = n9114 ^ n7081 ;
  assign n9155 = ~n9119 & ~n9154 ;
  assign n9156 = n9155 ^ n7081 ;
  assign n9157 = n9156 ^ n7383 ;
  assign n9151 = n9150 ^ n7542 ;
  assign n9152 = n8434 & n9151 ;
  assign n9153 = n9152 ^ n7542 ;
  assign n9158 = n9157 ^ n9153 ;
  assign n9160 = n9158 ^ x471 ;
  assign n9159 = n9158 ^ n9120 ;
  assign n9161 = n9160 ^ n9159 ;
  assign n9162 = n9125 & ~n9161 ;
  assign n9163 = n9162 ^ n9160 ;
  assign n9164 = n9163 ^ x470 ;
  assign n9145 = ~n9103 & n9126 ;
  assign n9165 = n9164 ^ n9145 ;
  assign n9140 = n9127 ^ n9101 ;
  assign n9141 = n9127 ^ n8546 ;
  assign n9142 = ~n9140 & n9141 ;
  assign n9143 = n9142 ^ n8546 ;
  assign n9144 = n9143 ^ n8586 ;
  assign n9166 = n9165 ^ n9144 ;
  assign n9167 = n8626 & n9166 ;
  assign n9168 = n9167 ^ n8016 ;
  assign n9135 = n9130 ^ n9099 ;
  assign n9136 = n9130 ^ n7595 ;
  assign n9137 = n9135 & ~n9136 ;
  assign n9138 = n9137 ^ n7595 ;
  assign n9139 = n9138 ^ n7592 ;
  assign n9169 = n9168 ^ n9139 ;
  assign n9170 = n9169 ^ x486 ;
  assign n9171 = n9170 ^ n9131 ;
  assign n9172 = n9171 ^ n9169 ;
  assign n9173 = n9134 & ~n9172 ;
  assign n9174 = n9173 ^ n9170 ;
  assign n9188 = n9156 ^ n9153 ;
  assign n9189 = n8453 ^ n7677 ;
  assign n9196 = n9195 ^ n9194 ;
  assign n9197 = ~n9189 & n9196 ;
  assign n9198 = n9197 ^ n7677 ;
  assign n9199 = n9198 ^ n7383 ;
  assign n9200 = n9199 ^ n9153 ;
  assign n9201 = n9200 ^ n9198 ;
  assign n9202 = ~n9188 & n9201 ;
  assign n9203 = n9202 ^ n9199 ;
  assign n9204 = n9203 ^ n7115 ;
  assign n9206 = n9204 ^ x470 ;
  assign n9205 = n9204 ^ n9158 ;
  assign n9207 = n9206 ^ n9205 ;
  assign n9208 = n9163 & ~n9207 ;
  assign n9209 = n9208 ^ n9206 ;
  assign n9210 = n9209 ^ x469 ;
  assign n9187 = ~n9145 & ~n9164 ;
  assign n9211 = n9210 ^ n9187 ;
  assign n9182 = n9165 ^ n9143 ;
  assign n9183 = n9165 ^ n8586 ;
  assign n9184 = ~n9182 & n9183 ;
  assign n9185 = n9184 ^ n8586 ;
  assign n9186 = n9185 ^ n8631 ;
  assign n9212 = n9211 ^ n9186 ;
  assign n9213 = n8648 & ~n9212 ;
  assign n9214 = n9213 ^ n8063 ;
  assign n9177 = n9168 ^ n9138 ;
  assign n9178 = n9168 ^ n7592 ;
  assign n9179 = ~n9177 & n9178 ;
  assign n9180 = n9179 ^ n7592 ;
  assign n9181 = n9180 ^ n7589 ;
  assign n9215 = n9214 ^ n9181 ;
  assign n9217 = n9215 ^ x485 ;
  assign n9216 = n9215 ^ n9169 ;
  assign n9218 = n9217 ^ n9216 ;
  assign n9219 = ~n9174 & n9218 ;
  assign n9220 = n9219 ^ n9217 ;
  assign n9238 = n8479 ^ n7686 ;
  assign n9245 = n9244 ^ n9243 ;
  assign n9246 = ~n9238 & n9245 ;
  assign n9247 = n9246 ^ n7686 ;
  assign n9234 = n9198 ^ n7115 ;
  assign n9235 = n9203 & ~n9234 ;
  assign n9236 = n9235 ^ n7115 ;
  assign n9237 = n9236 ^ n7130 ;
  assign n9248 = n9247 ^ n9237 ;
  assign n9250 = n9248 ^ x469 ;
  assign n9249 = n9248 ^ n9204 ;
  assign n9251 = n9250 ^ n9249 ;
  assign n9252 = ~n9209 & n9251 ;
  assign n9253 = n9252 ^ n9250 ;
  assign n9254 = n9253 ^ x468 ;
  assign n9233 = n9187 & n9210 ;
  assign n9255 = n9254 ^ n9233 ;
  assign n9228 = n9211 ^ n9185 ;
  assign n9229 = n9211 ^ n8631 ;
  assign n9230 = ~n9228 & ~n9229 ;
  assign n9231 = n9230 ^ n8631 ;
  assign n9232 = n9231 ^ n8676 ;
  assign n9256 = n9255 ^ n9232 ;
  assign n9257 = n8714 & n9256 ;
  assign n9258 = n9257 ^ n8107 ;
  assign n9223 = n9214 ^ n9180 ;
  assign n9224 = n9214 ^ n7589 ;
  assign n9225 = n9223 & n9224 ;
  assign n9226 = n9225 ^ n7589 ;
  assign n9227 = n9226 ^ n7585 ;
  assign n9259 = n9258 ^ n9227 ;
  assign n9261 = n9259 ^ x484 ;
  assign n9260 = n9259 ^ n9215 ;
  assign n9262 = n9261 ^ n9260 ;
  assign n9263 = ~n9220 & n9262 ;
  assign n9264 = n9263 ^ n9261 ;
  assign n9265 = n9264 ^ x483 ;
  assign n9096 = n9095 ^ x487 ;
  assign n9098 = n9097 ^ x486 ;
  assign n9132 = n9131 ^ n9098 ;
  assign n9133 = n9096 & ~n9132 ;
  assign n9175 = n9174 ^ x485 ;
  assign n9176 = n9133 & n9175 ;
  assign n9221 = n9220 ^ x484 ;
  assign n9222 = n9176 & n9221 ;
  assign n10621 = n9265 ^ n9222 ;
  assign n10069 = n8862 ^ n8819 ;
  assign n9837 = n8515 ^ x455 ;
  assign n9873 = n9837 ^ n9196 ;
  assign n9283 = n8501 ^ n7694 ;
  assign n9290 = n9289 ^ n9288 ;
  assign n9291 = n9283 & ~n9290 ;
  assign n9292 = n9291 ^ n7694 ;
  assign n9278 = n9247 ^ n9236 ;
  assign n9279 = n9247 ^ n7130 ;
  assign n9280 = ~n9278 & n9279 ;
  assign n9281 = n9280 ^ n7130 ;
  assign n9282 = n9281 ^ n7145 ;
  assign n9293 = n9292 ^ n9282 ;
  assign n9295 = n9293 ^ x468 ;
  assign n9294 = n9293 ^ n9248 ;
  assign n9296 = n9295 ^ n9294 ;
  assign n9297 = n9253 & ~n9296 ;
  assign n9298 = n9297 ^ n9295 ;
  assign n9328 = n8535 ^ n7703 ;
  assign n9335 = n9334 ^ n9333 ;
  assign n9336 = n9328 & n9335 ;
  assign n9337 = n9336 ^ n7703 ;
  assign n9323 = n9292 ^ n9281 ;
  assign n9324 = n9292 ^ n7145 ;
  assign n9325 = ~n9323 & ~n9324 ;
  assign n9326 = n9325 ^ n7145 ;
  assign n9327 = n9326 ^ n7156 ;
  assign n9338 = n9337 ^ n9327 ;
  assign n9340 = n9338 ^ x467 ;
  assign n9339 = n9338 ^ n9293 ;
  assign n9341 = n9340 ^ n9339 ;
  assign n9342 = ~n9298 & n9341 ;
  assign n9343 = n9342 ^ n9340 ;
  assign n9373 = n8575 ^ n7711 ;
  assign n9380 = n9379 ^ n9378 ;
  assign n9381 = ~n9373 & ~n9380 ;
  assign n9382 = n9381 ^ n7711 ;
  assign n9368 = n9337 ^ n9326 ;
  assign n9369 = n9337 ^ n7156 ;
  assign n9370 = ~n9368 & n9369 ;
  assign n9371 = n9370 ^ n7156 ;
  assign n9372 = n9371 ^ n7175 ;
  assign n9383 = n9382 ^ n9372 ;
  assign n9385 = n9383 ^ x466 ;
  assign n9384 = n9383 ^ n9338 ;
  assign n9386 = n9385 ^ n9384 ;
  assign n9387 = ~n9343 & n9386 ;
  assign n9388 = n9387 ^ n9385 ;
  assign n9418 = n8615 ^ n7539 ;
  assign n9425 = n9424 ^ n9423 ;
  assign n9426 = ~n9418 & ~n9425 ;
  assign n9427 = n9426 ^ n7539 ;
  assign n9413 = n9382 ^ n9371 ;
  assign n9414 = n9382 ^ n7175 ;
  assign n9415 = ~n9413 & ~n9414 ;
  assign n9416 = n9415 ^ n7175 ;
  assign n9417 = n9416 ^ n6869 ;
  assign n9428 = n9427 ^ n9417 ;
  assign n9430 = n9428 ^ x465 ;
  assign n9429 = n9428 ^ n9383 ;
  assign n9431 = n9430 ^ n9429 ;
  assign n9432 = n9388 & ~n9431 ;
  assign n9433 = n9432 ^ n9430 ;
  assign n9474 = n9428 ^ x464 ;
  assign n9475 = n9433 & ~n9474 ;
  assign n9476 = n9475 ^ x464 ;
  assign n9462 = n8660 ^ n7724 ;
  assign n9469 = n9468 ^ n9467 ;
  assign n9470 = n9462 & n9469 ;
  assign n9471 = n9470 ^ n7724 ;
  assign n9472 = n9471 ^ n7206 ;
  assign n9458 = n9427 ^ n9416 ;
  assign n9459 = n9427 ^ n6869 ;
  assign n9460 = n9458 & n9459 ;
  assign n9461 = n9460 ^ n6869 ;
  assign n9473 = n9472 ^ n9461 ;
  assign n9477 = n9476 ^ n9473 ;
  assign n9510 = n9471 ^ n9461 ;
  assign n9511 = ~n9472 & n9510 ;
  assign n9512 = n9511 ^ n7206 ;
  assign n9513 = n9512 ^ n7876 ;
  assign n9507 = n9506 ^ n7883 ;
  assign n9508 = ~n8702 & ~n9507 ;
  assign n9509 = n9508 ^ n7883 ;
  assign n9514 = n9513 ^ n9509 ;
  assign n9515 = n9514 ^ x479 ;
  assign n9516 = n9515 ^ n9476 ;
  assign n9517 = n9516 ^ n9514 ;
  assign n9518 = n9477 & n9517 ;
  assign n9519 = n9518 ^ n9515 ;
  assign n9549 = n8752 ^ n7962 ;
  assign n9557 = ~n9549 & ~n9556 ;
  assign n9558 = n9557 ^ n7962 ;
  assign n9545 = n9512 ^ n9509 ;
  assign n9546 = ~n9513 & ~n9545 ;
  assign n9547 = n9546 ^ n7876 ;
  assign n9548 = n9547 ^ n7246 ;
  assign n9559 = n9558 ^ n9548 ;
  assign n9561 = n9559 ^ x478 ;
  assign n9560 = n9559 ^ n9514 ;
  assign n9562 = n9561 ^ n9560 ;
  assign n9563 = n9519 & ~n9562 ;
  assign n9564 = n9563 ^ n9561 ;
  assign n9592 = n8794 ^ n8000 ;
  assign n9598 = n8399 ^ n8379 ;
  assign n9594 = n8794 ^ n8752 ;
  assign n9593 = n9555 ^ n8794 ;
  assign n9595 = n9594 ^ n9593 ;
  assign n9596 = ~n9554 & n9595 ;
  assign n9597 = n9596 ^ n9594 ;
  assign n9599 = n9598 ^ n9597 ;
  assign n9600 = n9592 & n9599 ;
  assign n9601 = n9600 ^ n8000 ;
  assign n9587 = n9558 ^ n9547 ;
  assign n9588 = n9558 ^ n7246 ;
  assign n9589 = ~n9587 & ~n9588 ;
  assign n9590 = n9589 ^ n7246 ;
  assign n9591 = n9590 ^ n7267 ;
  assign n9602 = n9601 ^ n9591 ;
  assign n9604 = n9602 ^ x477 ;
  assign n9603 = n9602 ^ n9559 ;
  assign n9605 = n9604 ^ n9603 ;
  assign n9606 = ~n9564 & n9605 ;
  assign n9607 = n9606 ^ n9604 ;
  assign n9636 = n8842 ^ n8051 ;
  assign n9642 = n8422 ^ n8400 ;
  assign n9638 = n8842 ^ n8794 ;
  assign n9637 = n9598 ^ n8842 ;
  assign n9639 = n9638 ^ n9637 ;
  assign n9640 = ~n9597 & n9639 ;
  assign n9641 = n9640 ^ n9638 ;
  assign n9643 = n9642 ^ n9641 ;
  assign n9644 = ~n9636 & ~n9643 ;
  assign n9645 = n9644 ^ n8051 ;
  assign n9631 = n9601 ^ n9590 ;
  assign n9632 = n9601 ^ n7267 ;
  assign n9633 = n9631 & n9632 ;
  assign n9634 = n9633 ^ n7267 ;
  assign n9635 = n9634 ^ n7291 ;
  assign n9646 = n9645 ^ n9635 ;
  assign n9648 = n9646 ^ x476 ;
  assign n9647 = n9646 ^ n9602 ;
  assign n9649 = n9648 ^ n9647 ;
  assign n9650 = ~n9607 & n9649 ;
  assign n9651 = n9650 ^ n9648 ;
  assign n9669 = n8883 ^ n8090 ;
  assign n9670 = n8444 ^ n8423 ;
  assign n9672 = n9670 ^ n8842 ;
  assign n9671 = n9670 ^ n9642 ;
  assign n9673 = n9672 ^ n9671 ;
  assign n9674 = n9641 & n9673 ;
  assign n9675 = n9674 ^ n9672 ;
  assign n9676 = n9675 ^ n8883 ;
  assign n9677 = ~n9669 & n9676 ;
  assign n9678 = n9677 ^ n8090 ;
  assign n9664 = n9645 ^ n9634 ;
  assign n9665 = n9645 ^ n7291 ;
  assign n9666 = n9664 & n9665 ;
  assign n9667 = n9666 ^ n7291 ;
  assign n9668 = n9667 ^ n7312 ;
  assign n9679 = n9678 ^ n9668 ;
  assign n9681 = n9679 ^ x475 ;
  assign n9680 = n9679 ^ n9646 ;
  assign n9682 = n9681 ^ n9680 ;
  assign n9683 = n9651 & ~n9682 ;
  assign n9684 = n9683 ^ n9681 ;
  assign n9723 = n8934 ^ n8139 ;
  assign n9729 = n8467 ^ n8445 ;
  assign n9725 = n8934 ^ n8883 ;
  assign n9724 = n9670 ^ n8934 ;
  assign n9726 = n9725 ^ n9724 ;
  assign n9727 = n9675 & ~n9726 ;
  assign n9728 = n9727 ^ n9725 ;
  assign n9730 = n9729 ^ n9728 ;
  assign n9731 = ~n9723 & ~n9730 ;
  assign n9732 = n9731 ^ n8139 ;
  assign n9718 = n9678 ^ n9667 ;
  assign n9719 = n9678 ^ n7312 ;
  assign n9720 = ~n9718 & ~n9719 ;
  assign n9721 = n9720 ^ n7312 ;
  assign n9722 = n9721 ^ n7490 ;
  assign n9733 = n9732 ^ n9722 ;
  assign n9735 = n9733 ^ x474 ;
  assign n9734 = n9733 ^ n9679 ;
  assign n9736 = n9735 ^ n9734 ;
  assign n9737 = n9684 & ~n9736 ;
  assign n9738 = n9737 ^ n9735 ;
  assign n9739 = n9738 ^ x473 ;
  assign n9685 = n9684 ^ x474 ;
  assign n9277 = ~n9233 & n9254 ;
  assign n9299 = n9298 ^ x467 ;
  assign n9322 = n9277 & ~n9299 ;
  assign n9344 = n9343 ^ x466 ;
  assign n9367 = n9322 & ~n9344 ;
  assign n9389 = n9388 ^ x465 ;
  assign n9412 = n9367 & n9389 ;
  assign n9434 = n9433 ^ x464 ;
  assign n9457 = ~n9412 & ~n9434 ;
  assign n9478 = n9477 ^ x479 ;
  assign n9501 = n9457 & ~n9478 ;
  assign n9520 = n9519 ^ x478 ;
  assign n9544 = ~n9501 & n9520 ;
  assign n9565 = n9564 ^ x477 ;
  assign n9586 = n9544 & ~n9565 ;
  assign n9608 = n9607 ^ x476 ;
  assign n9630 = ~n9586 & n9608 ;
  assign n9652 = n9651 ^ x475 ;
  assign n9686 = n9630 & ~n9652 ;
  assign n9717 = n9685 & ~n9686 ;
  assign n9740 = n9739 ^ n9717 ;
  assign n9653 = n9652 ^ n9630 ;
  assign n9609 = n9608 ^ n9586 ;
  assign n9566 = n9565 ^ n9544 ;
  assign n9521 = n9520 ^ n9501 ;
  assign n9479 = n9478 ^ n9457 ;
  assign n9435 = n9434 ^ n9412 ;
  assign n9390 = n9389 ^ n9367 ;
  assign n9345 = n9344 ^ n9322 ;
  assign n9300 = n9299 ^ n9277 ;
  assign n9272 = n9255 ^ n9231 ;
  assign n9273 = n9255 ^ n8676 ;
  assign n9274 = n9272 & ~n9273 ;
  assign n9275 = n9274 ^ n8676 ;
  assign n9317 = n9300 ^ n9275 ;
  assign n9318 = n9300 ^ n8719 ;
  assign n9319 = n9317 & ~n9318 ;
  assign n9320 = n9319 ^ n8719 ;
  assign n9362 = n9345 ^ n9320 ;
  assign n9363 = n9345 ^ n8764 ;
  assign n9364 = n9362 & n9363 ;
  assign n9365 = n9364 ^ n8764 ;
  assign n9407 = n9390 ^ n9365 ;
  assign n9408 = n9390 ^ n8809 ;
  assign n9409 = n9407 & ~n9408 ;
  assign n9410 = n9409 ^ n8809 ;
  assign n9452 = n9435 ^ n9410 ;
  assign n9453 = n9435 ^ n8853 ;
  assign n9454 = ~n9452 & ~n9453 ;
  assign n9455 = n9454 ^ n8853 ;
  assign n9496 = n9479 ^ n9455 ;
  assign n9497 = n9479 ^ n8899 ;
  assign n9498 = ~n9496 & n9497 ;
  assign n9499 = n9498 ^ n8899 ;
  assign n9539 = n9521 ^ n9499 ;
  assign n9540 = n9521 ^ n8945 ;
  assign n9541 = n9539 & n9540 ;
  assign n9542 = n9541 ^ n8945 ;
  assign n9581 = n9566 ^ n9542 ;
  assign n9582 = n9566 ^ n8988 ;
  assign n9583 = ~n9581 & n9582 ;
  assign n9584 = n9583 ^ n8988 ;
  assign n9625 = n9609 ^ n9584 ;
  assign n9626 = n9609 ^ n9005 ;
  assign n9627 = n9625 & ~n9626 ;
  assign n9628 = n9627 ^ n9005 ;
  assign n9688 = n9653 ^ n9628 ;
  assign n9689 = n9653 ^ n9029 ;
  assign n9690 = n9688 & ~n9689 ;
  assign n9691 = n9690 ^ n9029 ;
  assign n9687 = n9686 ^ n9685 ;
  assign n9712 = n9691 ^ n9687 ;
  assign n9713 = n9687 ^ n9057 ;
  assign n9714 = ~n9712 & ~n9713 ;
  assign n9715 = n9714 ^ n9057 ;
  assign n9817 = n9740 ^ n9715 ;
  assign n9818 = n9740 ^ n9074 ;
  assign n9819 = ~n9817 & n9818 ;
  assign n9820 = n9819 ^ n9074 ;
  assign n9812 = n7490 ^ x472 ;
  assign n9813 = n9812 ^ n8973 ;
  assign n9809 = n9732 ^ n9721 ;
  assign n9810 = n9732 ^ n7490 ;
  assign n9811 = n9809 & ~n9810 ;
  assign n9814 = n9813 ^ n9811 ;
  assign n9801 = n8979 ^ n8187 ;
  assign n9805 = n9729 ^ n8934 ;
  assign n9806 = ~n9728 & n9805 ;
  assign n9802 = n8488 ^ n8468 ;
  assign n9803 = n9802 ^ n8979 ;
  assign n9804 = n9803 ^ n9729 ;
  assign n9807 = n9806 ^ n9804 ;
  assign n9808 = ~n9801 & n9807 ;
  assign n9815 = n9814 ^ n9808 ;
  assign n9796 = n9733 ^ n9717 ;
  assign n9799 = ~n9738 & n9796 ;
  assign n9795 = n9738 ^ n9733 ;
  assign n9797 = n9796 ^ n9795 ;
  assign n9798 = ~x473 & ~n9797 ;
  assign n9800 = n9799 ^ n9798 ;
  assign n9816 = n9815 ^ n9800 ;
  assign n9838 = n9820 ^ n9816 ;
  assign n9839 = n9816 ^ n9111 ;
  assign n9840 = n9838 & n9839 ;
  assign n9841 = n9840 ^ n9111 ;
  assign n9842 = n9841 ^ n9837 ;
  assign n9870 = n9190 ^ n9150 ;
  assign n9871 = n9870 ^ n9837 ;
  assign n9872 = ~n9842 & n9871 ;
  assign n9874 = n9873 ^ n9872 ;
  assign n9947 = n9245 ^ n9196 ;
  assign n9946 = n9245 ^ n8550 ;
  assign n9948 = n9947 ^ n9946 ;
  assign n9949 = n9874 & n9948 ;
  assign n9950 = n9949 ^ n9946 ;
  assign n9967 = n8640 ^ n8596 ;
  assign n9969 = n9967 ^ n9245 ;
  assign n9951 = n8595 ^ n8550 ;
  assign n9968 = n9967 ^ n9951 ;
  assign n9970 = n9969 ^ n9968 ;
  assign n9971 = n9950 & ~n9970 ;
  assign n9972 = n9971 ^ n9969 ;
  assign n9989 = n9335 ^ n9290 ;
  assign n9988 = n9967 ^ n9335 ;
  assign n9990 = n9989 ^ n9988 ;
  assign n9991 = ~n9972 & ~n9990 ;
  assign n9992 = n9991 ^ n9989 ;
  assign n9993 = n8685 ^ n8641 ;
  assign n10010 = n9993 ^ n9335 ;
  assign n10011 = ~n9992 & n10010 ;
  assign n10012 = n10011 ^ n9335 ;
  assign n10009 = n8728 ^ n8686 ;
  assign n10013 = n10012 ^ n10009 ;
  assign n10030 = n9425 ^ n9380 ;
  assign n10029 = n10012 ^ n9425 ;
  assign n10031 = n10030 ^ n10029 ;
  assign n10032 = ~n10013 & ~n10031 ;
  assign n10033 = n10032 ^ n10030 ;
  assign n10034 = n8773 ^ n8729 ;
  assign n10047 = n10034 ^ n9425 ;
  assign n10048 = n10033 & ~n10047 ;
  assign n10049 = n10048 ^ n9425 ;
  assign n10045 = n8818 ^ n8774 ;
  assign n10065 = n10049 ^ n10045 ;
  assign n10066 = n10049 ^ n9469 ;
  assign n10067 = n10065 & ~n10066 ;
  assign n10068 = n10067 ^ n9469 ;
  assign n10070 = n10069 ^ n10068 ;
  assign n9939 = n9506 ^ n8703 ;
  assign n10616 = n10070 ^ n9939 ;
  assign n10091 = n8908 ^ n8863 ;
  assign n10087 = n10069 ^ n9939 ;
  assign n10088 = n10068 ^ n9939 ;
  assign n10089 = n10087 & n10088 ;
  assign n10086 = n10069 ^ n9556 ;
  assign n10090 = n10089 ^ n10086 ;
  assign n10092 = n10091 ^ n10090 ;
  assign n10619 = n10616 ^ n10092 ;
  assign n10046 = n10045 ^ n9469 ;
  assign n10050 = n10049 ^ n10046 ;
  assign n10035 = n10034 ^ n10033 ;
  assign n10313 = n10050 ^ n10035 ;
  assign n10223 = n9807 ^ n8979 ;
  assign n10112 = n9599 ^ n9556 ;
  assign n10111 = n10091 ^ n9599 ;
  assign n10113 = n10112 ^ n10111 ;
  assign n10114 = n10090 & ~n10113 ;
  assign n10115 = n10114 ^ n10112 ;
  assign n10133 = n9643 ^ n9599 ;
  assign n10116 = n8954 ^ n8909 ;
  assign n10132 = n10116 ^ n9643 ;
  assign n10134 = n10133 ^ n10132 ;
  assign n10135 = ~n10115 & ~n10134 ;
  assign n10136 = n10135 ^ n10133 ;
  assign n10153 = n9676 ^ n9643 ;
  assign n10137 = n8997 ^ n8955 ;
  assign n10152 = n10137 ^ n9676 ;
  assign n10154 = n10153 ^ n10152 ;
  assign n10155 = ~n10136 & ~n10154 ;
  assign n10156 = n10155 ^ n10153 ;
  assign n10174 = n9730 ^ n9676 ;
  assign n10157 = n9019 ^ n8998 ;
  assign n10173 = n10157 ^ n9730 ;
  assign n10175 = n10174 ^ n10173 ;
  assign n10176 = ~n10156 & ~n10175 ;
  assign n10177 = n10176 ^ n10174 ;
  assign n10178 = n9043 ^ n9020 ;
  assign n10227 = n10178 ^ n9730 ;
  assign n10228 = n10177 & n10227 ;
  assign n10225 = n9066 ^ n9044 ;
  assign n10224 = n10178 ^ n9807 ;
  assign n10226 = n10225 ^ n10224 ;
  assign n10229 = n10228 ^ n10226 ;
  assign n10230 = ~n10223 & ~n10229 ;
  assign n10220 = n8139 ^ x504 ;
  assign n10221 = n10220 ^ n9801 ;
  assign n10172 = n9730 ^ n8934 ;
  assign n10179 = n10178 ^ n10177 ;
  assign n10180 = n10172 & n10179 ;
  assign n10181 = n10180 ^ n8934 ;
  assign n10158 = n10157 ^ n10156 ;
  assign n10159 = ~n9675 & n10158 ;
  assign n10160 = n10159 ^ n8883 ;
  assign n10131 = n9643 ^ n8842 ;
  assign n10138 = n10137 ^ n10136 ;
  assign n10139 = n10131 & ~n10138 ;
  assign n10140 = n10139 ^ n8842 ;
  assign n10110 = n9599 ^ n8794 ;
  assign n10117 = n10116 ^ n10115 ;
  assign n10118 = ~n10110 & n10117 ;
  assign n10119 = n10118 ^ n8794 ;
  assign n10028 = n9425 ^ n8615 ;
  assign n10036 = n10028 & n10035 ;
  assign n10037 = n10036 ^ n8615 ;
  assign n10008 = n9380 ^ n8575 ;
  assign n10014 = n10013 ^ n9380 ;
  assign n10015 = n10008 & ~n10014 ;
  assign n10016 = n10015 ^ n8575 ;
  assign n9987 = n9335 ^ n8535 ;
  assign n9994 = n9993 ^ n9992 ;
  assign n9995 = n9987 & ~n9994 ;
  assign n9996 = n9995 ^ n8535 ;
  assign n9966 = n9290 ^ n8501 ;
  assign n9973 = n9972 ^ n9290 ;
  assign n9974 = n9966 & ~n9973 ;
  assign n9975 = n9974 ^ n8501 ;
  assign n9945 = n9245 ^ n8479 ;
  assign n9952 = n9951 ^ n9950 ;
  assign n9953 = n9945 & ~n9952 ;
  assign n9954 = n9953 ^ n8479 ;
  assign n9869 = n9196 ^ n8453 ;
  assign n9875 = n9874 ^ n8550 ;
  assign n9876 = ~n9869 & ~n9875 ;
  assign n9877 = n9876 ^ n8453 ;
  assign n9794 = n9111 ^ n8408 ;
  assign n9821 = n9820 ^ n9111 ;
  assign n9822 = n9821 ^ n9816 ;
  assign n9823 = ~n9794 & ~n9822 ;
  assign n9824 = n9823 ^ n8408 ;
  assign n9716 = n9715 ^ n9074 ;
  assign n9741 = n9740 ^ n9716 ;
  assign n9742 = ~n9073 & ~n9741 ;
  assign n9743 = n9742 ^ n8390 ;
  assign n9624 = n9029 ^ n8346 ;
  assign n9629 = n9628 ^ n9029 ;
  assign n9654 = n9653 ^ n9629 ;
  assign n9655 = n9624 & ~n9654 ;
  assign n9656 = n9655 ^ n8346 ;
  assign n9585 = n9584 ^ n9005 ;
  assign n9610 = n9609 ^ n9585 ;
  assign n9611 = ~n9022 & ~n9610 ;
  assign n9612 = n9611 ^ n8324 ;
  assign n9543 = n9542 ^ n8988 ;
  assign n9567 = n9566 ^ n9543 ;
  assign n9568 = ~n9001 & n9567 ;
  assign n9569 = n9568 ^ n8298 ;
  assign n9500 = n9499 ^ n8945 ;
  assign n9522 = n9521 ^ n9500 ;
  assign n9523 = n8983 & ~n9522 ;
  assign n9524 = n9523 ^ n8280 ;
  assign n9456 = n9455 ^ n8899 ;
  assign n9480 = n9479 ^ n9456 ;
  assign n9481 = ~n8917 & ~n9480 ;
  assign n9482 = n9481 ^ n8258 ;
  assign n9411 = n9410 ^ n8853 ;
  assign n9436 = n9435 ^ n9411 ;
  assign n9437 = n8894 & ~n9436 ;
  assign n9438 = n9437 ^ n8235 ;
  assign n9366 = n9365 ^ n8809 ;
  assign n9391 = n9390 ^ n9366 ;
  assign n9392 = n8825 & ~n9391 ;
  assign n9393 = n9392 ^ n8215 ;
  assign n9321 = n9320 ^ n8764 ;
  assign n9346 = n9345 ^ n9321 ;
  assign n9347 = n8805 & ~n9346 ;
  assign n9348 = n9347 ^ n8192 ;
  assign n9276 = n9275 ^ n8719 ;
  assign n9301 = n9300 ^ n9276 ;
  assign n9302 = ~n8736 & n9301 ;
  assign n9303 = n9302 ^ n8150 ;
  assign n9267 = n9258 ^ n9226 ;
  assign n9268 = n9258 ^ n7585 ;
  assign n9269 = ~n9267 & n9268 ;
  assign n9270 = n9269 ^ n7585 ;
  assign n9312 = n9303 ^ n9270 ;
  assign n9313 = n9303 ^ n7582 ;
  assign n9314 = n9312 & ~n9313 ;
  assign n9315 = n9314 ^ n7582 ;
  assign n9357 = n9348 ^ n9315 ;
  assign n9358 = n9348 ^ n7578 ;
  assign n9359 = n9357 & ~n9358 ;
  assign n9360 = n9359 ^ n7578 ;
  assign n9402 = n9393 ^ n9360 ;
  assign n9403 = n9393 ^ n7575 ;
  assign n9404 = n9402 & ~n9403 ;
  assign n9405 = n9404 ^ n7575 ;
  assign n9447 = n9438 ^ n9405 ;
  assign n9448 = n9438 ^ n7572 ;
  assign n9449 = ~n9447 & ~n9448 ;
  assign n9450 = n9449 ^ n7572 ;
  assign n9491 = n9482 ^ n9450 ;
  assign n9492 = n9482 ^ n7568 ;
  assign n9493 = ~n9491 & ~n9492 ;
  assign n9494 = n9493 ^ n7568 ;
  assign n9534 = n9524 ^ n9494 ;
  assign n9535 = n9524 ^ n7564 ;
  assign n9536 = n9534 & n9535 ;
  assign n9537 = n9536 ^ n7564 ;
  assign n9576 = n9569 ^ n9537 ;
  assign n9577 = n9569 ^ n7561 ;
  assign n9578 = n9576 & ~n9577 ;
  assign n9579 = n9578 ^ n7561 ;
  assign n9619 = n9612 ^ n9579 ;
  assign n9620 = n9612 ^ n7557 ;
  assign n9621 = n9619 & ~n9620 ;
  assign n9622 = n9621 ^ n7557 ;
  assign n9696 = n9656 ^ n9622 ;
  assign n9697 = n9656 ^ n7554 ;
  assign n9698 = ~n9696 & ~n9697 ;
  assign n9699 = n9698 ^ n7554 ;
  assign n9663 = n9057 ^ n8364 ;
  assign n9692 = n9691 ^ n9057 ;
  assign n9693 = n9692 ^ n9687 ;
  assign n9694 = n9663 & ~n9693 ;
  assign n9695 = n9694 ^ n8364 ;
  assign n9707 = n9699 ^ n9695 ;
  assign n9708 = n9695 ^ n7550 ;
  assign n9709 = ~n9707 & ~n9708 ;
  assign n9710 = n9709 ^ n7550 ;
  assign n9790 = n9743 ^ n9710 ;
  assign n9791 = n9743 ^ n7547 ;
  assign n9792 = ~n9790 & n9791 ;
  assign n9793 = n9792 ^ n7547 ;
  assign n9836 = n9824 ^ n9793 ;
  assign n9843 = n9842 ^ n9190 ;
  assign n9844 = n9150 & ~n9843 ;
  assign n9845 = n9844 ^ n9190 ;
  assign n9846 = n9845 ^ n7660 ;
  assign n9847 = n9846 ^ n9845 ;
  assign n9848 = n9847 ^ n9793 ;
  assign n9849 = n9836 & n9848 ;
  assign n9850 = n9849 ^ n9846 ;
  assign n9865 = n9845 ^ n7542 ;
  assign n9866 = n9850 & n9865 ;
  assign n9867 = n9866 ^ n7542 ;
  assign n9940 = n9877 ^ n9867 ;
  assign n9941 = n9877 ^ n7677 ;
  assign n9942 = ~n9940 & ~n9941 ;
  assign n9943 = n9942 ^ n7677 ;
  assign n9961 = n9954 ^ n9943 ;
  assign n9962 = n9954 ^ n7686 ;
  assign n9963 = ~n9961 & ~n9962 ;
  assign n9964 = n9963 ^ n7686 ;
  assign n9982 = n9975 ^ n9964 ;
  assign n9983 = n9975 ^ n7694 ;
  assign n9984 = ~n9982 & n9983 ;
  assign n9985 = n9984 ^ n7694 ;
  assign n10003 = n9996 ^ n9985 ;
  assign n10004 = n9996 ^ n7703 ;
  assign n10005 = n10003 & n10004 ;
  assign n10006 = n10005 ^ n7703 ;
  assign n10023 = n10016 ^ n10006 ;
  assign n10024 = n10016 ^ n7711 ;
  assign n10025 = n10023 & ~n10024 ;
  assign n10026 = n10025 ^ n7711 ;
  assign n10044 = n10037 ^ n10026 ;
  assign n10051 = n9469 ^ n8660 ;
  assign n10052 = ~n10050 & ~n10051 ;
  assign n10053 = n10052 ^ n8660 ;
  assign n10054 = n10053 ^ n7539 ;
  assign n10055 = n10054 ^ n10053 ;
  assign n10056 = n10055 ^ n10026 ;
  assign n10057 = n10044 & n10056 ;
  assign n10058 = n10057 ^ n10054 ;
  assign n10071 = n10070 ^ n8703 ;
  assign n10072 = n9506 & ~n10071 ;
  assign n10073 = n10072 ^ n8703 ;
  assign n10075 = n10073 ^ n7724 ;
  assign n10074 = n10073 ^ n10053 ;
  assign n10076 = n10075 ^ n10074 ;
  assign n10077 = n10058 & n10076 ;
  assign n10078 = n10077 ^ n10075 ;
  assign n10085 = n9556 ^ n8752 ;
  assign n10093 = ~n10085 & n10092 ;
  assign n10094 = n10093 ^ n8752 ;
  assign n10096 = n10094 ^ n7883 ;
  assign n10095 = n10094 ^ n10073 ;
  assign n10097 = n10096 ^ n10095 ;
  assign n10098 = ~n10078 & ~n10097 ;
  assign n10099 = n10098 ^ n10096 ;
  assign n10106 = n10094 ^ n7962 ;
  assign n10107 = ~n10099 & ~n10106 ;
  assign n10108 = n10107 ^ n7962 ;
  assign n10126 = n10119 ^ n10108 ;
  assign n10127 = n10119 ^ n8000 ;
  assign n10128 = ~n10126 & n10127 ;
  assign n10129 = n10128 ^ n8000 ;
  assign n10147 = n10140 ^ n10129 ;
  assign n10148 = n10140 ^ n8051 ;
  assign n10149 = ~n10147 & ~n10148 ;
  assign n10150 = n10149 ^ n8051 ;
  assign n10167 = n10160 ^ n10150 ;
  assign n10168 = n10160 ^ n8090 ;
  assign n10169 = n10167 & ~n10168 ;
  assign n10170 = n10169 ^ n8090 ;
  assign n10217 = n10181 ^ n10170 ;
  assign n10218 = n10181 ^ n8139 ;
  assign n10219 = n10217 & ~n10218 ;
  assign n10222 = n10221 ^ n10219 ;
  assign n10231 = n10230 ^ n10222 ;
  assign n9825 = n9824 ^ n7660 ;
  assign n9826 = n9825 ^ n9793 ;
  assign n9271 = n9270 ^ n7582 ;
  assign n9304 = n9303 ^ n9271 ;
  assign n9306 = n9304 ^ x483 ;
  assign n9305 = n9304 ^ n9259 ;
  assign n9307 = n9306 ^ n9305 ;
  assign n9308 = n9264 & ~n9307 ;
  assign n9309 = n9308 ^ n9306 ;
  assign n9316 = n9315 ^ n7578 ;
  assign n9349 = n9348 ^ n9316 ;
  assign n9351 = n9349 ^ x482 ;
  assign n9350 = n9349 ^ n9304 ;
  assign n9352 = n9351 ^ n9350 ;
  assign n9353 = ~n9309 & n9352 ;
  assign n9354 = n9353 ^ n9351 ;
  assign n9361 = n9360 ^ n7575 ;
  assign n9394 = n9393 ^ n9361 ;
  assign n9396 = n9394 ^ x481 ;
  assign n9395 = n9394 ^ n9349 ;
  assign n9397 = n9396 ^ n9395 ;
  assign n9398 = ~n9354 & n9397 ;
  assign n9399 = n9398 ^ n9396 ;
  assign n9406 = n9405 ^ n7572 ;
  assign n9439 = n9438 ^ n9406 ;
  assign n9441 = n9439 ^ x480 ;
  assign n9440 = n9439 ^ n9394 ;
  assign n9442 = n9441 ^ n9440 ;
  assign n9443 = ~n9399 & n9442 ;
  assign n9444 = n9443 ^ n9441 ;
  assign n9451 = n9450 ^ n7568 ;
  assign n9483 = n9482 ^ n9451 ;
  assign n9485 = n9483 ^ x495 ;
  assign n9484 = n9483 ^ n9439 ;
  assign n9486 = n9485 ^ n9484 ;
  assign n9487 = ~n9444 & n9486 ;
  assign n9488 = n9487 ^ n9485 ;
  assign n9495 = n9494 ^ n7564 ;
  assign n9525 = n9524 ^ n9495 ;
  assign n9527 = n9525 ^ x494 ;
  assign n9526 = n9525 ^ n9483 ;
  assign n9528 = n9527 ^ n9526 ;
  assign n9529 = n9488 & ~n9528 ;
  assign n9530 = n9529 ^ n9527 ;
  assign n9538 = n9537 ^ n7561 ;
  assign n9570 = n9569 ^ n9538 ;
  assign n9572 = n9570 ^ x493 ;
  assign n9571 = n9570 ^ n9525 ;
  assign n9573 = n9572 ^ n9571 ;
  assign n9574 = n9530 & ~n9573 ;
  assign n9575 = n9574 ^ n9572 ;
  assign n9580 = n9579 ^ n7557 ;
  assign n9613 = n9612 ^ n9580 ;
  assign n9615 = n9613 ^ x492 ;
  assign n9614 = n9613 ^ n9570 ;
  assign n9616 = n9615 ^ n9614 ;
  assign n9617 = n9575 & ~n9616 ;
  assign n9618 = n9617 ^ n9615 ;
  assign n9623 = n9622 ^ n7554 ;
  assign n9657 = n9656 ^ n9623 ;
  assign n9659 = n9657 ^ x491 ;
  assign n9658 = n9657 ^ n9613 ;
  assign n9660 = n9659 ^ n9658 ;
  assign n9661 = n9618 & ~n9660 ;
  assign n9662 = n9661 ^ n9659 ;
  assign n9700 = n9699 ^ n7550 ;
  assign n9701 = n9700 ^ n9695 ;
  assign n9703 = n9701 ^ x490 ;
  assign n9702 = n9701 ^ n9657 ;
  assign n9704 = n9703 ^ n9702 ;
  assign n9705 = n9662 & ~n9704 ;
  assign n9706 = n9705 ^ n9703 ;
  assign n9711 = n9710 ^ n7547 ;
  assign n9744 = n9743 ^ n9711 ;
  assign n9746 = n9744 ^ x489 ;
  assign n9745 = n9744 ^ n9701 ;
  assign n9747 = n9746 ^ n9745 ;
  assign n9748 = ~n9706 & n9747 ;
  assign n9749 = n9748 ^ n9746 ;
  assign n9786 = n9744 ^ x488 ;
  assign n9787 = ~n9749 & n9786 ;
  assign n9788 = n9787 ^ x488 ;
  assign n9835 = n9826 ^ n9788 ;
  assign n9851 = n9850 ^ n7542 ;
  assign n9852 = n9851 ^ x503 ;
  assign n9853 = n9852 ^ n9826 ;
  assign n9854 = n9853 ^ n9851 ;
  assign n9855 = n9835 & ~n9854 ;
  assign n9856 = n9855 ^ n9852 ;
  assign n9868 = n9867 ^ n7677 ;
  assign n9878 = n9877 ^ n9868 ;
  assign n9880 = n9878 ^ x502 ;
  assign n9879 = n9878 ^ n9851 ;
  assign n9881 = n9880 ^ n9879 ;
  assign n9882 = ~n9856 & n9881 ;
  assign n9883 = n9882 ^ n9880 ;
  assign n9944 = n9943 ^ n7686 ;
  assign n9955 = n9954 ^ n9944 ;
  assign n9957 = n9955 ^ x501 ;
  assign n9956 = n9955 ^ n9878 ;
  assign n9958 = n9957 ^ n9956 ;
  assign n9959 = ~n9883 & n9958 ;
  assign n9960 = n9959 ^ n9957 ;
  assign n9965 = n9964 ^ n7694 ;
  assign n9976 = n9975 ^ n9965 ;
  assign n9978 = n9976 ^ x500 ;
  assign n9977 = n9976 ^ n9955 ;
  assign n9979 = n9978 ^ n9977 ;
  assign n9980 = n9960 & ~n9979 ;
  assign n9981 = n9980 ^ n9978 ;
  assign n9986 = n9985 ^ n7703 ;
  assign n9997 = n9996 ^ n9986 ;
  assign n9999 = n9997 ^ x499 ;
  assign n9998 = n9997 ^ n9976 ;
  assign n10000 = n9999 ^ n9998 ;
  assign n10001 = n9981 & ~n10000 ;
  assign n10002 = n10001 ^ n9999 ;
  assign n10007 = n10006 ^ n7711 ;
  assign n10017 = n10016 ^ n10007 ;
  assign n10019 = n10017 ^ x498 ;
  assign n10018 = n10017 ^ n9997 ;
  assign n10020 = n10019 ^ n10018 ;
  assign n10021 = n10002 & ~n10020 ;
  assign n10022 = n10021 ^ n10019 ;
  assign n10027 = n10026 ^ n7539 ;
  assign n10038 = n10037 ^ n10027 ;
  assign n10040 = n10038 ^ x497 ;
  assign n10039 = n10038 ^ n10017 ;
  assign n10041 = n10040 ^ n10039 ;
  assign n10042 = n10022 & ~n10041 ;
  assign n10043 = n10042 ^ n10040 ;
  assign n10059 = n10058 ^ n7724 ;
  assign n10061 = n10059 ^ x496 ;
  assign n10060 = n10059 ^ n10038 ;
  assign n10062 = n10061 ^ n10060 ;
  assign n10063 = n10043 & ~n10062 ;
  assign n10064 = n10063 ^ n10061 ;
  assign n10079 = n10078 ^ n7883 ;
  assign n10081 = n10079 ^ x511 ;
  assign n10080 = n10079 ^ n10059 ;
  assign n10082 = n10081 ^ n10080 ;
  assign n10083 = ~n10064 & n10082 ;
  assign n10084 = n10083 ^ n10081 ;
  assign n10100 = n10099 ^ n7962 ;
  assign n10102 = n10100 ^ x510 ;
  assign n10101 = n10100 ^ n10079 ;
  assign n10103 = n10102 ^ n10101 ;
  assign n10104 = ~n10084 & n10103 ;
  assign n10105 = n10104 ^ n10102 ;
  assign n10109 = n10108 ^ n8000 ;
  assign n10120 = n10119 ^ n10109 ;
  assign n10122 = n10120 ^ x509 ;
  assign n10121 = n10120 ^ n10100 ;
  assign n10123 = n10122 ^ n10121 ;
  assign n10124 = n10105 & ~n10123 ;
  assign n10125 = n10124 ^ n10122 ;
  assign n10130 = n10129 ^ n8051 ;
  assign n10141 = n10140 ^ n10130 ;
  assign n10143 = n10141 ^ x508 ;
  assign n10142 = n10141 ^ n10120 ;
  assign n10144 = n10143 ^ n10142 ;
  assign n10145 = n10125 & ~n10144 ;
  assign n10146 = n10145 ^ n10143 ;
  assign n10151 = n10150 ^ n8090 ;
  assign n10161 = n10160 ^ n10151 ;
  assign n10163 = n10161 ^ x507 ;
  assign n10162 = n10161 ^ n10141 ;
  assign n10164 = n10163 ^ n10162 ;
  assign n10165 = ~n10146 & n10164 ;
  assign n10166 = n10165 ^ n10163 ;
  assign n10171 = n10170 ^ n8139 ;
  assign n10182 = n10181 ^ n10171 ;
  assign n10184 = n10182 ^ x506 ;
  assign n10183 = n10182 ^ n10161 ;
  assign n10185 = n10184 ^ n10183 ;
  assign n10186 = n10166 & ~n10185 ;
  assign n10187 = n10186 ^ n10184 ;
  assign n10189 = n10105 ^ x509 ;
  assign n9857 = n9856 ^ x502 ;
  assign n9789 = n9788 ^ x503 ;
  assign n9827 = n9826 ^ n9789 ;
  assign n9750 = n9749 ^ x488 ;
  assign n9751 = n9662 ^ x490 ;
  assign n9752 = n9618 ^ x491 ;
  assign n9753 = n9575 ^ x492 ;
  assign n9266 = n9222 & ~n9265 ;
  assign n9310 = n9309 ^ x482 ;
  assign n9311 = ~n9266 & ~n9310 ;
  assign n9355 = n9354 ^ x481 ;
  assign n9356 = ~n9311 & n9355 ;
  assign n9400 = n9399 ^ x480 ;
  assign n9401 = n9356 & n9400 ;
  assign n9445 = n9444 ^ x495 ;
  assign n9446 = n9401 & n9445 ;
  assign n9489 = n9488 ^ x494 ;
  assign n9490 = n9446 & ~n9489 ;
  assign n9531 = n9530 ^ x493 ;
  assign n9754 = n9490 & ~n9531 ;
  assign n9755 = n9753 & ~n9754 ;
  assign n9756 = ~n9752 & ~n9755 ;
  assign n9757 = ~n9751 & n9756 ;
  assign n9758 = n9706 ^ x489 ;
  assign n9759 = n9757 & n9758 ;
  assign n9828 = n9750 & n9759 ;
  assign n9858 = ~n9827 & n9828 ;
  assign n9864 = n9857 & n9858 ;
  assign n9884 = n9883 ^ x501 ;
  assign n10190 = ~n9864 & ~n9884 ;
  assign n10191 = n9960 ^ x500 ;
  assign n10192 = ~n10190 & ~n10191 ;
  assign n10193 = n9981 ^ x499 ;
  assign n10194 = ~n10192 & n10193 ;
  assign n10195 = n10002 ^ x498 ;
  assign n10196 = n10194 & n10195 ;
  assign n10197 = n10022 ^ x497 ;
  assign n10198 = ~n10196 & ~n10197 ;
  assign n10199 = n10043 ^ x496 ;
  assign n10200 = ~n10198 & n10199 ;
  assign n10201 = n10064 ^ x511 ;
  assign n10202 = n10200 & ~n10201 ;
  assign n10203 = n10084 ^ x510 ;
  assign n10204 = ~n10202 & n10203 ;
  assign n10205 = ~n10189 & n10204 ;
  assign n10206 = n10125 ^ x508 ;
  assign n10207 = ~n10205 & n10206 ;
  assign n10208 = n10146 ^ x507 ;
  assign n10209 = ~n10207 & n10208 ;
  assign n10210 = n10166 ^ x506 ;
  assign n10211 = n10209 & ~n10210 ;
  assign n10212 = n10211 ^ n10182 ;
  assign n10215 = n10187 & n10212 ;
  assign n10188 = n10187 ^ n10182 ;
  assign n10213 = n10212 ^ n10188 ;
  assign n10214 = x505 & n10213 ;
  assign n10216 = n10215 ^ n10214 ;
  assign n10232 = n10231 ^ n10216 ;
  assign n10233 = n10232 ^ n9994 ;
  assign n10234 = n10187 ^ x505 ;
  assign n10235 = n10234 ^ n10211 ;
  assign n10236 = n10235 ^ n9973 ;
  assign n10237 = n10208 ^ n10207 ;
  assign n10238 = n10237 ^ n9875 ;
  assign n10241 = n9870 ^ n9842 ;
  assign n10239 = n10206 ^ n10205 ;
  assign n10242 = n10241 ^ n10239 ;
  assign n10282 = n10204 ^ n10189 ;
  assign n10273 = n10201 ^ n10200 ;
  assign n10268 = n10199 ^ n10198 ;
  assign n10263 = n10197 ^ n10196 ;
  assign n10254 = n10193 ^ n10192 ;
  assign n10249 = n10191 ^ n10190 ;
  assign n9885 = n9884 ^ n9864 ;
  assign n9829 = n9828 ^ n9827 ;
  assign n9777 = n9758 ^ n9757 ;
  assign n9772 = n9756 ^ n9751 ;
  assign n9767 = n9755 ^ n9752 ;
  assign n9762 = n9754 ^ n9753 ;
  assign n9532 = n9531 ^ n9490 ;
  assign n9761 = ~n9091 & ~n9532 ;
  assign n9763 = n9762 ^ n9761 ;
  assign n9764 = n9762 ^ n9128 ;
  assign n9765 = ~n9763 & n9764 ;
  assign n9766 = n9765 ^ n9128 ;
  assign n9768 = n9767 ^ n9766 ;
  assign n9769 = n9767 ^ n9166 ;
  assign n9770 = ~n9768 & n9769 ;
  assign n9771 = n9770 ^ n9166 ;
  assign n9773 = n9772 ^ n9771 ;
  assign n9774 = n9772 ^ n9212 ;
  assign n9775 = n9773 & n9774 ;
  assign n9776 = n9775 ^ n9212 ;
  assign n9778 = n9777 ^ n9776 ;
  assign n9779 = n9777 ^ n9256 ;
  assign n9780 = n9778 & n9779 ;
  assign n9781 = n9780 ^ n9256 ;
  assign n9760 = n9759 ^ n9750 ;
  assign n9782 = n9781 ^ n9760 ;
  assign n9783 = n9781 ^ n9301 ;
  assign n9784 = ~n9782 & n9783 ;
  assign n9785 = n9784 ^ n9301 ;
  assign n9830 = n9829 ^ n9785 ;
  assign n9831 = n9829 ^ n9346 ;
  assign n9832 = n9830 & n9831 ;
  assign n9833 = n9832 ^ n9346 ;
  assign n9834 = n9833 ^ n9391 ;
  assign n9859 = n9858 ^ n9857 ;
  assign n9860 = n9859 ^ n9833 ;
  assign n9861 = n9834 & n9860 ;
  assign n9862 = n9861 ^ n9391 ;
  assign n10245 = n9885 ^ n9862 ;
  assign n10246 = n9885 ^ n9436 ;
  assign n10247 = ~n10245 & n10246 ;
  assign n10248 = n10247 ^ n9436 ;
  assign n10250 = n10249 ^ n10248 ;
  assign n10251 = n10249 ^ n9480 ;
  assign n10252 = n10250 & ~n10251 ;
  assign n10253 = n10252 ^ n9480 ;
  assign n10255 = n10254 ^ n10253 ;
  assign n10256 = n10254 ^ n9522 ;
  assign n10257 = n10255 & ~n10256 ;
  assign n10258 = n10257 ^ n9522 ;
  assign n10244 = n10195 ^ n10194 ;
  assign n10259 = n10258 ^ n10244 ;
  assign n10260 = n10258 ^ n9567 ;
  assign n10261 = ~n10259 & ~n10260 ;
  assign n10262 = n10261 ^ n9567 ;
  assign n10264 = n10263 ^ n10262 ;
  assign n10265 = n10263 ^ n9610 ;
  assign n10266 = ~n10264 & ~n10265 ;
  assign n10267 = n10266 ^ n9610 ;
  assign n10269 = n10268 ^ n10267 ;
  assign n10270 = n10268 ^ n9654 ;
  assign n10271 = n10269 & ~n10270 ;
  assign n10272 = n10271 ^ n9654 ;
  assign n10274 = n10273 ^ n10272 ;
  assign n10275 = n10273 ^ n9693 ;
  assign n10276 = n10274 & ~n10275 ;
  assign n10277 = n10276 ^ n9693 ;
  assign n10243 = n10203 ^ n10202 ;
  assign n10278 = n10277 ^ n10243 ;
  assign n10279 = n10277 ^ n9741 ;
  assign n10280 = ~n10278 & n10279 ;
  assign n10281 = n10280 ^ n9741 ;
  assign n10283 = n10282 ^ n10281 ;
  assign n10284 = n10239 ^ n9822 ;
  assign n10285 = n10284 ^ n10239 ;
  assign n10286 = n10285 ^ n10281 ;
  assign n10287 = ~n10283 & n10286 ;
  assign n10288 = n10287 ^ n10284 ;
  assign n10289 = n10242 & ~n10288 ;
  assign n10240 = n10239 ^ n10237 ;
  assign n10290 = n10289 ^ n10240 ;
  assign n10291 = n10238 & n10290 ;
  assign n10292 = n10291 ^ n9875 ;
  assign n10293 = n10292 ^ n9952 ;
  assign n10294 = n10210 ^ n10209 ;
  assign n10295 = n10294 ^ n10292 ;
  assign n10296 = n10293 & ~n10295 ;
  assign n10297 = n10296 ^ n9952 ;
  assign n10298 = n10297 ^ n10235 ;
  assign n10299 = ~n10236 & n10298 ;
  assign n10300 = n10299 ^ n9973 ;
  assign n10301 = n10300 ^ n10232 ;
  assign n10302 = ~n10233 & n10301 ;
  assign n10303 = n10302 ^ n9994 ;
  assign n10304 = n10303 ^ n10014 ;
  assign n10305 = n10035 ^ n9096 ;
  assign n10306 = n10305 ^ n10035 ;
  assign n10307 = n10306 ^ n10303 ;
  assign n10308 = ~n10304 & n10307 ;
  assign n10309 = n10308 ^ n10305 ;
  assign n10310 = n9132 ^ n9096 ;
  assign n10311 = n10310 ^ n10035 ;
  assign n10312 = ~n10309 & ~n10311 ;
  assign n10314 = n10313 ^ n10312 ;
  assign n10316 = n9175 ^ n9133 ;
  assign n10315 = n9221 ^ n9176 ;
  assign n10317 = n10316 ^ n10315 ;
  assign n10318 = n10317 ^ n10050 ;
  assign n10319 = n10318 ^ n10315 ;
  assign n10320 = n10314 & ~n10319 ;
  assign n10321 = n10320 ^ n10317 ;
  assign n10617 = n10616 ^ n10315 ;
  assign n10618 = ~n10321 & n10617 ;
  assign n10620 = n10619 ^ n10618 ;
  assign n10622 = n10621 ^ n10620 ;
  assign n10623 = n10622 ^ n10092 ;
  assign n10624 = ~n9556 & ~n10623 ;
  assign n10625 = n10624 ^ n10092 ;
  assign n10324 = n10316 ^ n10314 ;
  assign n10325 = n10324 ^ n10050 ;
  assign n10326 = n9469 & n10325 ;
  assign n10327 = n10326 ^ n10050 ;
  assign n10328 = n10327 ^ n8660 ;
  assign n10450 = n10310 ^ n10309 ;
  assign n10451 = n10450 ^ n10035 ;
  assign n10452 = ~n9425 & n10451 ;
  assign n10453 = n10452 ^ n10035 ;
  assign n10443 = n10303 ^ n9096 ;
  assign n10444 = ~n9380 & ~n10443 ;
  assign n10445 = n10444 ^ n10013 ;
  assign n10329 = n9335 & ~n10301 ;
  assign n10330 = n10329 ^ n9994 ;
  assign n10331 = n10330 ^ n8535 ;
  assign n10332 = n9245 & n10295 ;
  assign n10333 = n10332 ^ n9952 ;
  assign n10334 = n10333 ^ n8479 ;
  assign n10335 = n9196 & ~n10290 ;
  assign n10336 = n10335 ^ n9875 ;
  assign n10337 = n10336 ^ n8453 ;
  assign n10338 = ~n9870 & n10288 ;
  assign n10339 = n10338 ^ n9842 ;
  assign n10340 = n10339 ^ n9190 ;
  assign n10343 = ~n9074 & n10278 ;
  assign n10344 = n10343 ^ n9741 ;
  assign n10345 = n10344 ^ n8390 ;
  assign n10410 = ~n9057 & ~n10274 ;
  assign n10411 = n10410 ^ n9693 ;
  assign n10404 = n9029 & ~n10269 ;
  assign n10405 = n10404 ^ n9654 ;
  assign n10398 = n9005 & n10264 ;
  assign n10399 = n10398 ^ n9610 ;
  assign n10392 = n8988 & n10259 ;
  assign n10393 = n10392 ^ n9567 ;
  assign n10386 = n8945 & ~n10255 ;
  assign n10387 = n10386 ^ n9522 ;
  assign n10380 = ~n8899 & ~n10250 ;
  assign n10381 = n10380 ^ n9480 ;
  assign n10374 = ~n8853 & n10245 ;
  assign n10375 = n10374 ^ n9436 ;
  assign n10368 = n8809 & ~n9860 ;
  assign n10369 = n10368 ^ n9391 ;
  assign n10362 = n8764 & ~n9830 ;
  assign n10363 = n10362 ^ n9346 ;
  assign n10356 = ~n8719 & n9782 ;
  assign n10357 = n10356 ^ n9301 ;
  assign n10350 = ~n8676 & ~n9778 ;
  assign n10351 = n10350 ^ n9256 ;
  assign n9919 = ~n8631 & ~n9773 ;
  assign n9920 = n9919 ^ n9212 ;
  assign n9904 = n8586 & n9768 ;
  assign n9905 = n9904 ^ n9166 ;
  assign n9894 = n8546 & n9763 ;
  assign n9895 = n9894 ^ n9128 ;
  assign n9887 = ~n9090 & n9532 ;
  assign n9888 = n9887 ^ n9089 ;
  assign n9892 = n8520 & n9888 ;
  assign n9899 = n9895 ^ n9892 ;
  assign n9900 = n9895 ^ n7977 ;
  assign n9901 = ~n9899 & ~n9900 ;
  assign n9902 = n9901 ^ n7977 ;
  assign n9914 = n9905 ^ n9902 ;
  assign n9915 = n9905 ^ n8016 ;
  assign n9916 = n9914 & n9915 ;
  assign n9917 = n9916 ^ n8016 ;
  assign n10346 = n9920 ^ n9917 ;
  assign n10347 = n9920 ^ n8063 ;
  assign n10348 = n10346 & n10347 ;
  assign n10349 = n10348 ^ n8063 ;
  assign n10352 = n10351 ^ n10349 ;
  assign n10353 = n10351 ^ n8107 ;
  assign n10354 = n10352 & ~n10353 ;
  assign n10355 = n10354 ^ n8107 ;
  assign n10358 = n10357 ^ n10355 ;
  assign n10359 = n10357 ^ n8150 ;
  assign n10360 = n10358 & n10359 ;
  assign n10361 = n10360 ^ n8150 ;
  assign n10364 = n10363 ^ n10361 ;
  assign n10365 = n10363 ^ n8192 ;
  assign n10366 = n10364 & ~n10365 ;
  assign n10367 = n10366 ^ n8192 ;
  assign n10370 = n10369 ^ n10367 ;
  assign n10371 = n10369 ^ n8215 ;
  assign n10372 = n10370 & ~n10371 ;
  assign n10373 = n10372 ^ n8215 ;
  assign n10376 = n10375 ^ n10373 ;
  assign n10377 = n10375 ^ n8235 ;
  assign n10378 = n10376 & n10377 ;
  assign n10379 = n10378 ^ n8235 ;
  assign n10382 = n10381 ^ n10379 ;
  assign n10383 = n10381 ^ n8258 ;
  assign n10384 = ~n10382 & ~n10383 ;
  assign n10385 = n10384 ^ n8258 ;
  assign n10388 = n10387 ^ n10385 ;
  assign n10389 = n10387 ^ n8280 ;
  assign n10390 = n10388 & ~n10389 ;
  assign n10391 = n10390 ^ n8280 ;
  assign n10394 = n10393 ^ n10391 ;
  assign n10395 = n10393 ^ n8298 ;
  assign n10396 = ~n10394 & ~n10395 ;
  assign n10397 = n10396 ^ n8298 ;
  assign n10400 = n10399 ^ n10397 ;
  assign n10401 = n10399 ^ n8324 ;
  assign n10402 = ~n10400 & n10401 ;
  assign n10403 = n10402 ^ n8324 ;
  assign n10406 = n10405 ^ n10403 ;
  assign n10407 = n10405 ^ n8346 ;
  assign n10408 = ~n10406 & ~n10407 ;
  assign n10409 = n10408 ^ n8346 ;
  assign n10412 = n10411 ^ n10409 ;
  assign n10413 = n10344 ^ n8364 ;
  assign n10414 = n10413 ^ n10344 ;
  assign n10415 = n10414 ^ n10409 ;
  assign n10416 = n10412 & ~n10415 ;
  assign n10417 = n10416 ^ n10413 ;
  assign n10418 = ~n10345 & ~n10417 ;
  assign n10419 = n10418 ^ n8390 ;
  assign n10341 = n9111 & n10283 ;
  assign n10342 = n10341 ^ n9822 ;
  assign n10420 = n10419 ^ n10342 ;
  assign n10421 = n10339 ^ n8408 ;
  assign n10422 = n10421 ^ n10339 ;
  assign n10423 = n10422 ^ n10342 ;
  assign n10424 = n10420 & n10423 ;
  assign n10425 = n10424 ^ n10421 ;
  assign n10426 = n10340 & ~n10425 ;
  assign n10427 = n10426 ^ n9190 ;
  assign n10428 = n10427 ^ n10336 ;
  assign n10429 = n10337 & ~n10428 ;
  assign n10430 = n10429 ^ n8453 ;
  assign n10431 = n10430 ^ n10333 ;
  assign n10432 = ~n10334 & ~n10431 ;
  assign n10433 = n10432 ^ n8479 ;
  assign n10434 = n10433 ^ n8501 ;
  assign n10435 = ~n9290 & n10298 ;
  assign n10436 = n10435 ^ n9972 ;
  assign n10437 = n10436 ^ n10433 ;
  assign n10438 = ~n10434 & ~n10437 ;
  assign n10439 = n10438 ^ n8501 ;
  assign n10440 = n10439 ^ n10330 ;
  assign n10441 = ~n10331 & ~n10440 ;
  assign n10442 = n10441 ^ n8535 ;
  assign n10446 = n10445 ^ n10442 ;
  assign n10447 = n10445 ^ n8575 ;
  assign n10448 = ~n10446 & ~n10447 ;
  assign n10449 = n10448 ^ n8575 ;
  assign n10454 = n10453 ^ n10449 ;
  assign n10455 = n10327 ^ n8615 ;
  assign n10456 = n10455 ^ n10327 ;
  assign n10457 = n10456 ^ n10449 ;
  assign n10458 = n10454 & n10457 ;
  assign n10459 = n10458 ^ n10455 ;
  assign n10460 = n10328 & ~n10459 ;
  assign n10461 = n10460 ^ n8660 ;
  assign n10462 = n10461 ^ n8703 ;
  assign n10322 = ~n9939 & ~n10321 ;
  assign n10323 = n10322 ^ n10070 ;
  assign n10612 = n10461 ^ n10323 ;
  assign n10613 = n10462 & ~n10612 ;
  assign n10614 = n10613 ^ n8703 ;
  assign n10615 = n10614 ^ n8752 ;
  assign n10626 = n10625 ^ n10615 ;
  assign n10463 = n10462 ^ n10323 ;
  assign n10464 = n10463 ^ x62 ;
  assign n10466 = n10449 ^ n8615 ;
  assign n10467 = n10466 ^ n10453 ;
  assign n10468 = n10467 ^ x48 ;
  assign n10471 = n10417 ^ n8390 ;
  assign n10472 = n10471 ^ x40 ;
  assign n10475 = n10355 ^ n8150 ;
  assign n10476 = n10475 ^ n10357 ;
  assign n10477 = n10476 ^ x34 ;
  assign n9893 = n9892 ^ n7977 ;
  assign n9896 = n9895 ^ n9893 ;
  assign n9889 = n9888 ^ n8520 ;
  assign n9890 = x39 & n9889 ;
  assign n9898 = n9896 ^ n9890 ;
  assign n9903 = n9902 ^ n8016 ;
  assign n9906 = n9905 ^ n9903 ;
  assign n9907 = n9906 ^ x38 ;
  assign n9908 = n9907 ^ n9896 ;
  assign n9909 = n9908 ^ n9906 ;
  assign n9910 = n9898 & ~n9909 ;
  assign n9911 = n9910 ^ n9907 ;
  assign n9918 = n9917 ^ n8063 ;
  assign n9921 = n9920 ^ n9918 ;
  assign n9923 = n9921 ^ x37 ;
  assign n9922 = n9921 ^ n9906 ;
  assign n9924 = n9923 ^ n9922 ;
  assign n9925 = n9911 & ~n9924 ;
  assign n9926 = n9925 ^ n9923 ;
  assign n10478 = n10349 ^ n8107 ;
  assign n10479 = n10478 ^ n10351 ;
  assign n10481 = n10479 ^ x36 ;
  assign n10480 = n10479 ^ n9921 ;
  assign n10482 = n10481 ^ n10480 ;
  assign n10483 = ~n9926 & n10482 ;
  assign n10484 = n10483 ^ n10481 ;
  assign n10486 = n10476 ^ x35 ;
  assign n10485 = n10479 ^ n10476 ;
  assign n10487 = n10486 ^ n10485 ;
  assign n10488 = ~n10484 & n10487 ;
  assign n10489 = n10488 ^ n10486 ;
  assign n10490 = ~n10477 & n10489 ;
  assign n10491 = n10490 ^ x34 ;
  assign n10473 = n10361 ^ n8192 ;
  assign n10474 = n10473 ^ n10363 ;
  assign n10492 = n10491 ^ n10474 ;
  assign n10493 = n10367 ^ n8215 ;
  assign n10494 = n10493 ^ n10369 ;
  assign n10495 = n10494 ^ x33 ;
  assign n10496 = n10495 ^ n10474 ;
  assign n10497 = n10496 ^ n10494 ;
  assign n10498 = n10492 & ~n10497 ;
  assign n10499 = n10498 ^ n10495 ;
  assign n10500 = n10373 ^ n8235 ;
  assign n10501 = n10500 ^ n10375 ;
  assign n10503 = n10501 ^ x32 ;
  assign n10502 = n10501 ^ n10494 ;
  assign n10504 = n10503 ^ n10502 ;
  assign n10505 = n10499 & ~n10504 ;
  assign n10506 = n10505 ^ n10503 ;
  assign n10507 = n10379 ^ n8258 ;
  assign n10508 = n10507 ^ n10381 ;
  assign n10510 = n10508 ^ x47 ;
  assign n10509 = n10508 ^ n10501 ;
  assign n10511 = n10510 ^ n10509 ;
  assign n10512 = ~n10506 & n10511 ;
  assign n10513 = n10512 ^ n10510 ;
  assign n10514 = n10385 ^ n8280 ;
  assign n10515 = n10514 ^ n10387 ;
  assign n10517 = n10515 ^ x46 ;
  assign n10516 = n10515 ^ n10508 ;
  assign n10518 = n10517 ^ n10516 ;
  assign n10519 = ~n10513 & n10518 ;
  assign n10520 = n10519 ^ n10517 ;
  assign n10521 = n10391 ^ n8298 ;
  assign n10522 = n10521 ^ n10393 ;
  assign n10524 = n10522 ^ x45 ;
  assign n10523 = n10522 ^ n10515 ;
  assign n10525 = n10524 ^ n10523 ;
  assign n10526 = n10520 & ~n10525 ;
  assign n10527 = n10526 ^ n10524 ;
  assign n10528 = n10397 ^ n8324 ;
  assign n10529 = n10528 ^ n10399 ;
  assign n10531 = n10529 ^ x44 ;
  assign n10530 = n10529 ^ n10522 ;
  assign n10532 = n10531 ^ n10530 ;
  assign n10533 = n10527 & ~n10532 ;
  assign n10534 = n10533 ^ n10531 ;
  assign n10535 = n10403 ^ n8346 ;
  assign n10536 = n10535 ^ n10405 ;
  assign n10538 = n10536 ^ x43 ;
  assign n10537 = n10536 ^ n10529 ;
  assign n10539 = n10538 ^ n10537 ;
  assign n10540 = n10534 & ~n10539 ;
  assign n10541 = n10540 ^ n10538 ;
  assign n10542 = n10409 ^ n8364 ;
  assign n10543 = n10542 ^ n10411 ;
  assign n10545 = n10543 ^ x42 ;
  assign n10544 = n10543 ^ n10536 ;
  assign n10546 = n10545 ^ n10544 ;
  assign n10547 = ~n10541 & n10546 ;
  assign n10548 = n10547 ^ n10545 ;
  assign n10550 = n10471 ^ x41 ;
  assign n10549 = n10543 ^ n10471 ;
  assign n10551 = n10550 ^ n10549 ;
  assign n10552 = ~n10548 & n10551 ;
  assign n10553 = n10552 ^ n10550 ;
  assign n10554 = n10472 & ~n10553 ;
  assign n10555 = n10554 ^ x40 ;
  assign n10469 = n10342 ^ n8408 ;
  assign n10470 = n10469 ^ n10419 ;
  assign n10556 = n10555 ^ n10470 ;
  assign n10557 = n10425 ^ n9190 ;
  assign n10558 = n10557 ^ x55 ;
  assign n10559 = n10558 ^ n10470 ;
  assign n10560 = n10559 ^ n10557 ;
  assign n10561 = ~n10556 & n10560 ;
  assign n10562 = n10561 ^ n10558 ;
  assign n10563 = n10427 ^ n8453 ;
  assign n10564 = n10563 ^ n10336 ;
  assign n10566 = n10564 ^ x54 ;
  assign n10565 = n10564 ^ n10557 ;
  assign n10567 = n10566 ^ n10565 ;
  assign n10568 = n10562 & ~n10567 ;
  assign n10569 = n10568 ^ n10566 ;
  assign n10570 = n10430 ^ n8479 ;
  assign n10571 = n10570 ^ n10333 ;
  assign n10573 = n10571 ^ x53 ;
  assign n10572 = n10571 ^ n10564 ;
  assign n10574 = n10573 ^ n10572 ;
  assign n10575 = n10569 & ~n10574 ;
  assign n10576 = n10575 ^ n10573 ;
  assign n10577 = n10436 ^ n10434 ;
  assign n10579 = n10577 ^ x52 ;
  assign n10578 = n10577 ^ n10571 ;
  assign n10580 = n10579 ^ n10578 ;
  assign n10581 = ~n10576 & n10580 ;
  assign n10582 = n10581 ^ n10579 ;
  assign n10583 = n10439 ^ n8535 ;
  assign n10584 = n10583 ^ n10330 ;
  assign n10586 = n10584 ^ x51 ;
  assign n10585 = n10584 ^ n10577 ;
  assign n10587 = n10586 ^ n10585 ;
  assign n10588 = n10582 & ~n10587 ;
  assign n10589 = n10588 ^ n10586 ;
  assign n10590 = n10442 ^ n8575 ;
  assign n10591 = n10590 ^ n10445 ;
  assign n10593 = n10591 ^ x50 ;
  assign n10592 = n10591 ^ n10584 ;
  assign n10594 = n10593 ^ n10592 ;
  assign n10595 = ~n10589 & n10594 ;
  assign n10596 = n10595 ^ n10593 ;
  assign n10598 = n10467 ^ x49 ;
  assign n10597 = n10591 ^ n10467 ;
  assign n10599 = n10598 ^ n10597 ;
  assign n10600 = n10596 & ~n10599 ;
  assign n10601 = n10600 ^ n10598 ;
  assign n10602 = n10468 & ~n10601 ;
  assign n10603 = n10602 ^ x48 ;
  assign n10465 = n10459 ^ n8660 ;
  assign n10604 = n10603 ^ n10465 ;
  assign n10607 = n10465 ^ x63 ;
  assign n10608 = n10604 & ~n10607 ;
  assign n10605 = n10463 ^ x63 ;
  assign n10609 = n10608 ^ n10605 ;
  assign n10610 = ~n10464 & n10609 ;
  assign n10611 = n10610 ^ x62 ;
  assign n10627 = n10626 ^ n10611 ;
  assign n10628 = n10625 ^ n10614 ;
  assign n10634 = n9310 ^ n9266 ;
  assign n10630 = n10117 ^ n10092 ;
  assign n10629 = n10621 ^ n10117 ;
  assign n10631 = n10630 ^ n10629 ;
  assign n10632 = ~n10620 & ~n10631 ;
  assign n10633 = n10632 ^ n10629 ;
  assign n10635 = n10634 ^ n10633 ;
  assign n10636 = n10635 ^ n10117 ;
  assign n10637 = n9599 & n10636 ;
  assign n10638 = n10637 ^ n10117 ;
  assign n10639 = n10638 ^ n8752 ;
  assign n10640 = n10639 ^ n10614 ;
  assign n10641 = n10640 ^ n10638 ;
  assign n10642 = n10628 & ~n10641 ;
  assign n10643 = n10642 ^ n10639 ;
  assign n10644 = n10643 ^ n8794 ;
  assign n10645 = n10644 ^ x61 ;
  assign n10646 = n10645 ^ n10611 ;
  assign n10647 = n10646 ^ n10644 ;
  assign n10648 = n10627 & n10647 ;
  assign n10649 = n10648 ^ n10645 ;
  assign n10762 = n10649 ^ x60 ;
  assign n10711 = n10527 ^ x44 ;
  assign n9891 = n9890 ^ x38 ;
  assign n9897 = n9896 ^ n9891 ;
  assign n9912 = n9911 ^ x37 ;
  assign n9913 = ~n9897 & ~n9912 ;
  assign n9927 = n9926 ^ x36 ;
  assign n10712 = n9913 & n9927 ;
  assign n10713 = n10484 ^ x35 ;
  assign n10714 = n10712 & n10713 ;
  assign n10715 = n10489 ^ x34 ;
  assign n10716 = ~n10714 & n10715 ;
  assign n10717 = n10491 ^ x33 ;
  assign n10718 = n10717 ^ n10474 ;
  assign n10719 = n10716 & n10718 ;
  assign n10720 = n10499 ^ x32 ;
  assign n10721 = ~n10719 & ~n10720 ;
  assign n10722 = n10506 ^ x47 ;
  assign n10723 = ~n10721 & ~n10722 ;
  assign n10724 = n10513 ^ x46 ;
  assign n10725 = ~n10723 & n10724 ;
  assign n10726 = n10520 ^ x45 ;
  assign n10727 = ~n10725 & n10726 ;
  assign n10728 = ~n10711 & ~n10727 ;
  assign n10729 = n10534 ^ x43 ;
  assign n10730 = n10728 & ~n10729 ;
  assign n10731 = n10541 ^ x42 ;
  assign n10732 = ~n10730 & ~n10731 ;
  assign n10733 = n10548 ^ x41 ;
  assign n10734 = ~n10732 & n10733 ;
  assign n10735 = n10553 ^ x40 ;
  assign n10736 = n10734 & n10735 ;
  assign n10737 = n10555 ^ x55 ;
  assign n10738 = n10737 ^ n10470 ;
  assign n10739 = n10736 & n10738 ;
  assign n10740 = n10562 ^ x54 ;
  assign n10741 = ~n10739 & n10740 ;
  assign n10742 = n10569 ^ x53 ;
  assign n10743 = n10741 & n10742 ;
  assign n10744 = n10576 ^ x52 ;
  assign n10745 = n10743 & ~n10744 ;
  assign n10746 = n10582 ^ x51 ;
  assign n10747 = n10745 & n10746 ;
  assign n10748 = n10589 ^ x50 ;
  assign n10749 = ~n10747 & n10748 ;
  assign n10750 = n10596 ^ x49 ;
  assign n10751 = n10749 & ~n10750 ;
  assign n10752 = n10601 ^ x48 ;
  assign n10753 = n10751 & n10752 ;
  assign n10754 = n10603 ^ x63 ;
  assign n10755 = n10754 ^ n10465 ;
  assign n10756 = n10753 & ~n10755 ;
  assign n10757 = n10609 ^ x62 ;
  assign n10758 = ~n10756 & n10757 ;
  assign n10759 = n10611 ^ x61 ;
  assign n10760 = n10759 ^ n10626 ;
  assign n10761 = n10758 & n10760 ;
  assign n10800 = n10762 ^ n10761 ;
  assign n10844 = ~n9091 & ~n10800 ;
  assign n10845 = n10844 ^ n9532 ;
  assign n10846 = ~n9090 & ~n10845 ;
  assign n10847 = n10846 ^ n8546 ;
  assign n10659 = n9355 ^ n9311 ;
  assign n10655 = n10138 ^ n10117 ;
  assign n10654 = n10634 ^ n10138 ;
  assign n10656 = n10655 ^ n10654 ;
  assign n10657 = ~n10633 & ~n10656 ;
  assign n10658 = n10657 ^ n10655 ;
  assign n10660 = n10659 ^ n10658 ;
  assign n10661 = n10660 ^ n10138 ;
  assign n10662 = ~n9643 & ~n10661 ;
  assign n10663 = n10662 ^ n10138 ;
  assign n10650 = n10638 ^ n8794 ;
  assign n10651 = ~n10643 & ~n10650 ;
  assign n10652 = n10651 ^ n8794 ;
  assign n10653 = n10652 ^ n8842 ;
  assign n10664 = n10663 ^ n10653 ;
  assign n10666 = n10664 ^ x60 ;
  assign n10665 = n10664 ^ n10644 ;
  assign n10667 = n10666 ^ n10665 ;
  assign n10668 = n10649 & ~n10667 ;
  assign n10669 = n10668 ^ n10666 ;
  assign n10764 = n10669 ^ x59 ;
  assign n10763 = ~n10761 & ~n10762 ;
  assign n10805 = n10764 ^ n10763 ;
  assign n9533 = n9532 ^ n9091 ;
  assign n10801 = n9533 & n10800 ;
  assign n10806 = n10805 ^ n10801 ;
  assign n10848 = n9128 & n10806 ;
  assign n10802 = n9761 ^ n9128 ;
  assign n10803 = n10802 ^ n9762 ;
  assign n10849 = n10848 ^ n10803 ;
  assign n10850 = n10849 ^ n10846 ;
  assign n10851 = n10847 & ~n10850 ;
  assign n10852 = n10851 ^ n8546 ;
  assign n10853 = n10852 ^ n8586 ;
  assign n10804 = n10803 ^ n10801 ;
  assign n10807 = n10804 & ~n10806 ;
  assign n10808 = n10807 ^ n10803 ;
  assign n10675 = n9400 ^ n9356 ;
  assign n10677 = n10675 ^ n10138 ;
  assign n10676 = n10675 ^ n10659 ;
  assign n10678 = n10677 ^ n10676 ;
  assign n10679 = ~n10658 & n10678 ;
  assign n10680 = n10679 ^ n10677 ;
  assign n10681 = n9676 & ~n10680 ;
  assign n10682 = n10681 ^ n10158 ;
  assign n10670 = n10663 ^ n10652 ;
  assign n10671 = n10663 ^ n8842 ;
  assign n10672 = ~n10670 & n10671 ;
  assign n10673 = n10672 ^ n8842 ;
  assign n10674 = n10673 ^ n8883 ;
  assign n10683 = n10682 ^ n10674 ;
  assign n10685 = n10683 ^ x59 ;
  assign n10684 = n10683 ^ n10664 ;
  assign n10686 = n10685 ^ n10684 ;
  assign n10687 = n10669 & ~n10686 ;
  assign n10688 = n10687 ^ n10685 ;
  assign n10766 = n10688 ^ x58 ;
  assign n10765 = ~n10763 & n10764 ;
  assign n10798 = n10766 ^ n10765 ;
  assign n10854 = n10808 ^ n10798 ;
  assign n10855 = n9166 & n10854 ;
  assign n10796 = n9766 ^ n9166 ;
  assign n10797 = n10796 ^ n9767 ;
  assign n10856 = n10855 ^ n10797 ;
  assign n10857 = n10856 ^ n10852 ;
  assign n10858 = n10853 & ~n10857 ;
  assign n10859 = n10858 ^ n8586 ;
  assign n10860 = n10859 ^ n8631 ;
  assign n10799 = n10798 ^ n10797 ;
  assign n10809 = n10808 ^ n10797 ;
  assign n10810 = n10799 & ~n10809 ;
  assign n10811 = n10810 ^ n10798 ;
  assign n10699 = n9445 ^ n9401 ;
  assign n10695 = n10179 ^ n10158 ;
  assign n10694 = n10675 ^ n10179 ;
  assign n10696 = n10695 ^ n10694 ;
  assign n10697 = n10680 & n10696 ;
  assign n10698 = n10697 ^ n10695 ;
  assign n10700 = n10699 ^ n10698 ;
  assign n10701 = n10700 ^ n10179 ;
  assign n10702 = ~n9730 & n10701 ;
  assign n10703 = n10702 ^ n10179 ;
  assign n10689 = n10682 ^ n10673 ;
  assign n10690 = n10682 ^ n8883 ;
  assign n10691 = n10689 & ~n10690 ;
  assign n10692 = n10691 ^ n8883 ;
  assign n10693 = n10692 ^ n8934 ;
  assign n10704 = n10703 ^ n10693 ;
  assign n10706 = n10704 ^ x58 ;
  assign n10705 = n10704 ^ n10683 ;
  assign n10707 = n10706 ^ n10705 ;
  assign n10708 = ~n10688 & n10707 ;
  assign n10709 = n10708 ^ n10706 ;
  assign n10791 = n10709 ^ x57 ;
  assign n10767 = n10765 & ~n10766 ;
  assign n10792 = n10791 ^ n10767 ;
  assign n10812 = n10811 ^ n10792 ;
  assign n10861 = ~n9212 & n10812 ;
  assign n10793 = n9771 ^ n9212 ;
  assign n10794 = n10793 ^ n9772 ;
  assign n10862 = n10861 ^ n10794 ;
  assign n10863 = n10862 ^ n10859 ;
  assign n10864 = ~n10860 & ~n10863 ;
  assign n10865 = n10864 ^ n8631 ;
  assign n10866 = n10865 ^ n8676 ;
  assign n10795 = n10794 ^ n10792 ;
  assign n10813 = n10795 & ~n10812 ;
  assign n10814 = n10813 ^ n10794 ;
  assign n10783 = n10699 ^ n10179 ;
  assign n10784 = ~n10698 & n10783 ;
  assign n10781 = n9489 ^ n9446 ;
  assign n10780 = n10699 ^ n10229 ;
  assign n10782 = n10781 ^ n10780 ;
  assign n10785 = n10784 ^ n10782 ;
  assign n10786 = n10785 ^ n10229 ;
  assign n10787 = n9807 & ~n10786 ;
  assign n10777 = n10229 ^ n8979 ;
  assign n10776 = n8934 ^ x56 ;
  assign n10778 = n10777 ^ n10776 ;
  assign n10773 = n10703 ^ n10692 ;
  assign n10774 = n10703 ^ n8934 ;
  assign n10775 = n10773 & ~n10774 ;
  assign n10779 = n10778 ^ n10775 ;
  assign n10788 = n10787 ^ n10779 ;
  assign n10768 = n10767 ^ n10704 ;
  assign n10771 = ~n10709 & n10768 ;
  assign n10710 = n10709 ^ n10704 ;
  assign n10769 = n10768 ^ n10710 ;
  assign n10770 = x57 & n10769 ;
  assign n10772 = n10771 ^ n10770 ;
  assign n10789 = n10788 ^ n10772 ;
  assign n10867 = n10814 ^ n10789 ;
  assign n10868 = n9256 & ~n10867 ;
  assign n9937 = n9776 ^ n9256 ;
  assign n9938 = n9937 ^ n9777 ;
  assign n10869 = n10868 ^ n9938 ;
  assign n10870 = n10869 ^ n10865 ;
  assign n10871 = n10866 & ~n10870 ;
  assign n10872 = n10871 ^ n8676 ;
  assign n9934 = n9783 ^ n9760 ;
  assign n10817 = n10789 ^ n9934 ;
  assign n10790 = n10789 ^ n9938 ;
  assign n10815 = n10814 ^ n9938 ;
  assign n10816 = n10790 & n10815 ;
  assign n10818 = n10817 ^ n10816 ;
  assign n9935 = n9889 ^ x39 ;
  assign n10840 = n10818 ^ n9935 ;
  assign n10841 = n10840 ^ n9934 ;
  assign n10842 = n9301 & ~n10841 ;
  assign n10843 = n10842 ^ n9934 ;
  assign n10873 = n10872 ^ n10843 ;
  assign n10874 = n10872 ^ n8719 ;
  assign n10875 = n10873 & n10874 ;
  assign n10876 = n10875 ^ n8719 ;
  assign n11011 = n10876 ^ n8764 ;
  assign n9936 = n9935 ^ n9934 ;
  assign n10819 = n9936 & n10818 ;
  assign n10820 = n10819 ^ n9935 ;
  assign n10877 = n10820 ^ n9897 ;
  assign n10878 = ~n9346 & n10877 ;
  assign n10821 = n9785 ^ n9346 ;
  assign n10822 = n10821 ^ n9829 ;
  assign n10879 = n10878 ^ n10822 ;
  assign n11012 = n11011 ^ n10879 ;
  assign n11013 = n11012 ^ x193 ;
  assign n11015 = n10845 ^ n9090 ;
  assign n11016 = x199 & n11015 ;
  assign n11014 = n10849 ^ n10847 ;
  assign n11017 = n11016 ^ n11014 ;
  assign n11018 = n10856 ^ n10853 ;
  assign n11019 = n11018 ^ x198 ;
  assign n11020 = n11019 ^ n11014 ;
  assign n11021 = n11020 ^ n11018 ;
  assign n11022 = ~n11017 & n11021 ;
  assign n11023 = n11022 ^ n11019 ;
  assign n11024 = n10862 ^ n10860 ;
  assign n11026 = n11024 ^ x197 ;
  assign n11025 = n11024 ^ n11018 ;
  assign n11027 = n11026 ^ n11025 ;
  assign n11028 = ~n11023 & n11027 ;
  assign n11029 = n11028 ^ n11026 ;
  assign n11030 = n10869 ^ n10866 ;
  assign n11032 = n11030 ^ x196 ;
  assign n11031 = n11030 ^ n11024 ;
  assign n11033 = n11032 ^ n11031 ;
  assign n11034 = n11029 & ~n11033 ;
  assign n11035 = n11034 ^ n11032 ;
  assign n11036 = n10874 ^ n10843 ;
  assign n11038 = n11036 ^ x195 ;
  assign n11037 = n11036 ^ n11030 ;
  assign n11039 = n11038 ^ n11037 ;
  assign n11040 = n11035 & ~n11039 ;
  assign n11041 = n11040 ^ n11038 ;
  assign n11043 = n11012 ^ x194 ;
  assign n11042 = n11036 ^ n11012 ;
  assign n11044 = n11043 ^ n11042 ;
  assign n11045 = ~n11041 & n11044 ;
  assign n11046 = n11045 ^ n11043 ;
  assign n11047 = ~n11013 & n11046 ;
  assign n11048 = n11047 ^ x193 ;
  assign n10823 = n10822 ^ n10820 ;
  assign n9930 = n9860 ^ n9391 ;
  assign n10824 = n9930 ^ n9897 ;
  assign n10825 = n10824 ^ n9930 ;
  assign n10826 = n10825 ^ n10820 ;
  assign n10827 = ~n10823 & n10826 ;
  assign n10828 = n10827 ^ n10824 ;
  assign n9932 = n9912 ^ n9897 ;
  assign n10885 = n10828 ^ n9932 ;
  assign n10886 = n10885 ^ n9860 ;
  assign n10887 = ~n9391 & ~n10886 ;
  assign n10888 = n10887 ^ n9860 ;
  assign n10880 = n10879 ^ n10876 ;
  assign n10881 = n10879 ^ n8764 ;
  assign n10882 = n10880 & n10881 ;
  assign n10883 = n10882 ^ n8764 ;
  assign n10884 = n10883 ^ n8809 ;
  assign n11010 = n10888 ^ n10884 ;
  assign n11049 = n11048 ^ n11010 ;
  assign n10889 = n10888 ^ n10883 ;
  assign n10890 = n10884 & n10889 ;
  assign n10891 = n10890 ^ n8809 ;
  assign n11050 = n10891 ^ n8853 ;
  assign n9933 = n9932 ^ n9930 ;
  assign n10829 = n9933 & n10828 ;
  assign n9863 = n9862 ^ n9436 ;
  assign n9886 = n9885 ^ n9863 ;
  assign n9931 = n9930 ^ n9886 ;
  assign n10830 = n10829 ^ n9931 ;
  assign n9928 = n9927 ^ n9913 ;
  assign n10892 = n10830 ^ n9928 ;
  assign n10893 = n10892 ^ n9886 ;
  assign n10894 = ~n9436 & n10893 ;
  assign n10895 = n10894 ^ n9886 ;
  assign n11051 = n11050 ^ n10895 ;
  assign n11052 = n11051 ^ x192 ;
  assign n11053 = n11052 ^ n11010 ;
  assign n11054 = n11053 ^ n11051 ;
  assign n11055 = n11049 & ~n11054 ;
  assign n11056 = n11055 ^ n11052 ;
  assign n10896 = n10895 ^ n10891 ;
  assign n10897 = n10895 ^ n8853 ;
  assign n10898 = n10896 & n10897 ;
  assign n10899 = n10898 ^ n8853 ;
  assign n11057 = n10899 ^ n8899 ;
  assign n10836 = n10248 ^ n9480 ;
  assign n10837 = n10836 ^ n10249 ;
  assign n10833 = n10713 ^ n10712 ;
  assign n9929 = n9928 ^ n9886 ;
  assign n10831 = ~n9929 & n10830 ;
  assign n10832 = n10831 ^ n9928 ;
  assign n10834 = n10833 ^ n10832 ;
  assign n10835 = ~n9480 & n10834 ;
  assign n10838 = n10837 ^ n10835 ;
  assign n11058 = n11057 ^ n10838 ;
  assign n11060 = n11058 ^ x207 ;
  assign n11059 = n11058 ^ n11051 ;
  assign n11061 = n11060 ^ n11059 ;
  assign n11062 = ~n11056 & n11061 ;
  assign n11063 = n11062 ^ n11060 ;
  assign n10839 = n10838 ^ n8899 ;
  assign n10900 = n10899 ^ n10838 ;
  assign n10901 = ~n10839 & n10900 ;
  assign n10902 = n10901 ^ n8899 ;
  assign n11064 = n10902 ^ n8945 ;
  assign n10906 = n10253 ^ n9522 ;
  assign n10907 = n10906 ^ n10254 ;
  assign n10908 = n10907 ^ n10837 ;
  assign n10904 = n10837 ^ n10832 ;
  assign n10905 = ~n10834 & n10904 ;
  assign n10909 = n10908 ^ n10905 ;
  assign n10903 = n10715 ^ n10714 ;
  assign n10910 = n10909 ^ n10903 ;
  assign n10911 = n10910 ^ n10907 ;
  assign n10912 = ~n9522 & n10911 ;
  assign n10913 = n10912 ^ n10907 ;
  assign n11065 = n11064 ^ n10913 ;
  assign n11067 = n11065 ^ x206 ;
  assign n11066 = n11065 ^ n11058 ;
  assign n11068 = n11067 ^ n11066 ;
  assign n11069 = ~n11063 & n11068 ;
  assign n11070 = n11069 ^ n11067 ;
  assign n11267 = n11070 ^ x205 ;
  assign n11259 = n11046 ^ x193 ;
  assign n11260 = n11010 ^ x192 ;
  assign n11261 = n11260 ^ n11048 ;
  assign n11262 = ~n11259 & ~n11261 ;
  assign n11263 = n11056 ^ x207 ;
  assign n11264 = ~n11262 & ~n11263 ;
  assign n11265 = n11063 ^ x206 ;
  assign n11266 = n11264 & ~n11265 ;
  assign n11585 = n11267 ^ n11266 ;
  assign n11571 = n11263 ^ n11262 ;
  assign n11002 = n10282 ^ n9822 ;
  assign n11003 = n11002 ^ n10281 ;
  assign n10918 = n10260 ^ n10244 ;
  assign n10919 = n10918 ^ n10907 ;
  assign n10920 = n10919 ^ n10918 ;
  assign n10921 = n10920 ^ n10903 ;
  assign n10922 = n10909 & n10921 ;
  assign n10923 = n10922 ^ n10919 ;
  assign n10933 = n10262 ^ n9610 ;
  assign n10934 = n10933 ^ n10263 ;
  assign n10936 = n10934 ^ n10918 ;
  assign n10924 = n10718 ^ n10716 ;
  assign n10935 = n10934 ^ n10924 ;
  assign n10937 = n10936 ^ n10935 ;
  assign n10938 = n10923 & ~n10937 ;
  assign n10939 = n10938 ^ n10936 ;
  assign n10949 = n10267 ^ n9654 ;
  assign n10950 = n10949 ^ n10268 ;
  assign n10952 = n10950 ^ n10934 ;
  assign n10940 = n10720 ^ n10719 ;
  assign n10951 = n10950 ^ n10940 ;
  assign n10953 = n10952 ^ n10951 ;
  assign n10954 = ~n10939 & ~n10953 ;
  assign n10955 = n10954 ^ n10952 ;
  assign n10965 = n10272 ^ n9693 ;
  assign n10966 = n10965 ^ n10273 ;
  assign n10968 = n10966 ^ n10950 ;
  assign n10956 = n10722 ^ n10721 ;
  assign n10967 = n10966 ^ n10956 ;
  assign n10969 = n10968 ^ n10967 ;
  assign n10970 = ~n10955 & ~n10969 ;
  assign n10971 = n10970 ^ n10968 ;
  assign n10981 = n10279 ^ n10243 ;
  assign n10983 = n10981 ^ n10966 ;
  assign n10972 = n10724 ^ n10723 ;
  assign n10982 = n10981 ^ n10972 ;
  assign n10984 = n10983 ^ n10982 ;
  assign n10985 = n10971 & ~n10984 ;
  assign n10986 = n10985 ^ n10983 ;
  assign n10987 = n10726 ^ n10725 ;
  assign n10997 = n10987 ^ n10981 ;
  assign n10998 = ~n10986 & ~n10997 ;
  assign n10999 = n10998 ^ n10981 ;
  assign n10996 = n10727 ^ n10711 ;
  assign n11000 = n10999 ^ n10996 ;
  assign n11559 = n11003 ^ n11000 ;
  assign n11558 = n11261 ^ n11259 ;
  assign n11560 = n11559 ^ n11558 ;
  assign n10988 = n10987 ^ n10986 ;
  assign n11562 = n11259 ^ n10988 ;
  assign n10925 = n10924 ^ n10923 ;
  assign n11535 = n10925 ^ n10910 ;
  assign n11300 = n11015 ^ x199 ;
  assign n11298 = n10837 ^ n10834 ;
  assign n11301 = n11300 ^ n11298 ;
  assign n11226 = n10740 ^ n10739 ;
  assign n11130 = n10290 ^ n9875 ;
  assign n11127 = n10288 ^ n10241 ;
  assign n11131 = n11130 ^ n11127 ;
  assign n11110 = n10729 ^ n10728 ;
  assign n11111 = n11110 ^ n10999 ;
  assign n11108 = n11003 ^ n10999 ;
  assign n11109 = ~n11000 & n11108 ;
  assign n11112 = n11111 ^ n11109 ;
  assign n11128 = n11127 ^ n11110 ;
  assign n11129 = ~n11112 & n11128 ;
  assign n11132 = n11131 ^ n11129 ;
  assign n11151 = n10294 ^ n10293 ;
  assign n11152 = n11151 ^ n11130 ;
  assign n11153 = n11152 ^ n11151 ;
  assign n11126 = n10731 ^ n10730 ;
  assign n11154 = n11153 ^ n11126 ;
  assign n11155 = ~n11132 & ~n11154 ;
  assign n11156 = n11155 ^ n11152 ;
  assign n11173 = n10297 ^ n9973 ;
  assign n11174 = n11173 ^ n10235 ;
  assign n11176 = n11174 ^ n11151 ;
  assign n11157 = n10733 ^ n10732 ;
  assign n11175 = n11174 ^ n11157 ;
  assign n11177 = n11176 ^ n11175 ;
  assign n11178 = ~n11156 & n11177 ;
  assign n11179 = n11178 ^ n11176 ;
  assign n11196 = n10300 ^ n9994 ;
  assign n11197 = n11196 ^ n10232 ;
  assign n11199 = n11197 ^ n11174 ;
  assign n11180 = n10735 ^ n10734 ;
  assign n11198 = n11197 ^ n11180 ;
  assign n11200 = n11199 ^ n11198 ;
  assign n11201 = ~n11179 & n11200 ;
  assign n11202 = n11201 ^ n11199 ;
  assign n11219 = n10014 ^ n9096 ;
  assign n11220 = n11219 ^ n10303 ;
  assign n11222 = n11220 ^ n11197 ;
  assign n11203 = n10738 ^ n10736 ;
  assign n11221 = n11220 ^ n11203 ;
  assign n11223 = n11222 ^ n11221 ;
  assign n11224 = n11202 & n11223 ;
  assign n11225 = n11224 ^ n11222 ;
  assign n11227 = n11226 ^ n11225 ;
  assign n11228 = n11227 ^ n11220 ;
  assign n11229 = ~n10014 & n11228 ;
  assign n11230 = n11229 ^ n11220 ;
  assign n11204 = n11203 ^ n11202 ;
  assign n11205 = n11204 ^ n11197 ;
  assign n11206 = ~n9994 & n11205 ;
  assign n11207 = n11206 ^ n11197 ;
  assign n11181 = n11180 ^ n11179 ;
  assign n11182 = n11181 ^ n11174 ;
  assign n11183 = ~n9973 & ~n11182 ;
  assign n11184 = n11183 ^ n11174 ;
  assign n11158 = n11157 ^ n11156 ;
  assign n11159 = n11158 ^ n11151 ;
  assign n11160 = ~n9952 & ~n11159 ;
  assign n11161 = n11160 ^ n11151 ;
  assign n11001 = ~n9822 & ~n11000 ;
  assign n11004 = n11003 ^ n11001 ;
  assign n10989 = n10988 ^ n10981 ;
  assign n10990 = ~n9741 & n10989 ;
  assign n10991 = n10990 ^ n10981 ;
  assign n10973 = n10972 ^ n10971 ;
  assign n10974 = n10973 ^ n10966 ;
  assign n10975 = ~n9693 & ~n10974 ;
  assign n10976 = n10975 ^ n10966 ;
  assign n10957 = n10956 ^ n10955 ;
  assign n10958 = n10957 ^ n10950 ;
  assign n10959 = ~n9654 & n10958 ;
  assign n10960 = n10959 ^ n10950 ;
  assign n10941 = n10940 ^ n10939 ;
  assign n10942 = n10941 ^ n10934 ;
  assign n10943 = ~n9610 & n10942 ;
  assign n10944 = n10943 ^ n10934 ;
  assign n10926 = n10925 ^ n10918 ;
  assign n10927 = n9567 & ~n10926 ;
  assign n10928 = n10927 ^ n10918 ;
  assign n10914 = n10913 ^ n10902 ;
  assign n10915 = n10913 ^ n8945 ;
  assign n10916 = n10914 & n10915 ;
  assign n10917 = n10916 ^ n8945 ;
  assign n10929 = n10928 ^ n10917 ;
  assign n10930 = n10928 ^ n8988 ;
  assign n10931 = ~n10929 & n10930 ;
  assign n10932 = n10931 ^ n8988 ;
  assign n10945 = n10944 ^ n10932 ;
  assign n10946 = n10944 ^ n9005 ;
  assign n10947 = n10945 & ~n10946 ;
  assign n10948 = n10947 ^ n9005 ;
  assign n10961 = n10960 ^ n10948 ;
  assign n10962 = n10960 ^ n9029 ;
  assign n10963 = ~n10961 & n10962 ;
  assign n10964 = n10963 ^ n9029 ;
  assign n10977 = n10976 ^ n10964 ;
  assign n10978 = n10976 ^ n9057 ;
  assign n10979 = ~n10977 & ~n10978 ;
  assign n10980 = n10979 ^ n9057 ;
  assign n10992 = n10991 ^ n10980 ;
  assign n10993 = n10991 ^ n9074 ;
  assign n10994 = ~n10992 & n10993 ;
  assign n10995 = n10994 ^ n9074 ;
  assign n11107 = n11004 ^ n10995 ;
  assign n11113 = n10241 & ~n11112 ;
  assign n11114 = n11113 ^ n10288 ;
  assign n11115 = n11114 ^ n9111 ;
  assign n11116 = n11115 ^ n11114 ;
  assign n11117 = n11116 ^ n10995 ;
  assign n11118 = ~n11107 & ~n11117 ;
  assign n11119 = n11118 ^ n11115 ;
  assign n11137 = n11114 ^ n9870 ;
  assign n11138 = n11119 & n11137 ;
  assign n11139 = n11138 ^ n9870 ;
  assign n11140 = n11139 ^ n9196 ;
  assign n11133 = n11132 ^ n11126 ;
  assign n11134 = n11133 ^ n10290 ;
  assign n11135 = ~n9875 & ~n11134 ;
  assign n11136 = n11135 ^ n10290 ;
  assign n11147 = n11139 ^ n11136 ;
  assign n11148 = ~n11140 & ~n11147 ;
  assign n11149 = n11148 ^ n9196 ;
  assign n11168 = n11161 ^ n11149 ;
  assign n11169 = n11161 ^ n9245 ;
  assign n11170 = n11168 & ~n11169 ;
  assign n11171 = n11170 ^ n9245 ;
  assign n11191 = n11184 ^ n11171 ;
  assign n11192 = n11184 ^ n9290 ;
  assign n11193 = ~n11191 & ~n11192 ;
  assign n11194 = n11193 ^ n9290 ;
  assign n11214 = n11207 ^ n11194 ;
  assign n11215 = n11207 ^ n9335 ;
  assign n11216 = n11214 & n11215 ;
  assign n11217 = n11216 ^ n9335 ;
  assign n11246 = n11230 ^ n11217 ;
  assign n11247 = n11230 ^ n9380 ;
  assign n11248 = n11246 & n11247 ;
  assign n11249 = n11248 ^ n9380 ;
  assign n11241 = n10742 ^ n10741 ;
  assign n11238 = n11226 ^ n11220 ;
  assign n11239 = ~n11225 & ~n11238 ;
  assign n11237 = n11220 ^ n10450 ;
  assign n11240 = n11239 ^ n11237 ;
  assign n11242 = n11241 ^ n11240 ;
  assign n11243 = n11242 ^ n10450 ;
  assign n11244 = n10035 & n11243 ;
  assign n11245 = n11244 ^ n10450 ;
  assign n11305 = n11249 ^ n11245 ;
  assign n11306 = n10744 ^ n10743 ;
  assign n11307 = n11306 ^ n10450 ;
  assign n11308 = n11307 ^ n11241 ;
  assign n11309 = n11308 ^ n11306 ;
  assign n11310 = ~n11240 & ~n11309 ;
  assign n11311 = n11310 ^ n11307 ;
  assign n11312 = ~n10050 & n11311 ;
  assign n11313 = n11312 ^ n10324 ;
  assign n11314 = n11313 ^ n9425 ;
  assign n11315 = n11314 ^ n11313 ;
  assign n11316 = n11315 ^ n11249 ;
  assign n11317 = n11305 & n11316 ;
  assign n11318 = n11317 ^ n11314 ;
  assign n11335 = n11313 ^ n9469 ;
  assign n11336 = ~n11318 & ~n11335 ;
  assign n11337 = n11336 ^ n9469 ;
  assign n11338 = n11337 ^ n9939 ;
  assign n11330 = n10746 ^ n10745 ;
  assign n11324 = n10616 ^ n10321 ;
  assign n11326 = n11324 ^ n10324 ;
  assign n11325 = n11324 ^ n11306 ;
  assign n11327 = n11326 ^ n11325 ;
  assign n11328 = ~n11311 & ~n11327 ;
  assign n11329 = n11328 ^ n11326 ;
  assign n11331 = n11330 ^ n11329 ;
  assign n11332 = n11331 ^ n10321 ;
  assign n11333 = ~n10616 & n11332 ;
  assign n11334 = n11333 ^ n11331 ;
  assign n11339 = n11338 ^ n11334 ;
  assign n11319 = n11318 ^ n9469 ;
  assign n11007 = n10980 ^ n9074 ;
  assign n11008 = n11007 ^ n10991 ;
  assign n11009 = n11008 ^ x200 ;
  assign n11071 = n10917 ^ n8988 ;
  assign n11072 = n11071 ^ n10928 ;
  assign n11074 = n11072 ^ x205 ;
  assign n11073 = n11072 ^ n11065 ;
  assign n11075 = n11074 ^ n11073 ;
  assign n11076 = n11070 & ~n11075 ;
  assign n11077 = n11076 ^ n11074 ;
  assign n11078 = n10932 ^ n9005 ;
  assign n11079 = n11078 ^ n10944 ;
  assign n11081 = n11079 ^ x204 ;
  assign n11080 = n11079 ^ n11072 ;
  assign n11082 = n11081 ^ n11080 ;
  assign n11083 = ~n11077 & n11082 ;
  assign n11084 = n11083 ^ n11081 ;
  assign n11085 = n10948 ^ n9029 ;
  assign n11086 = n11085 ^ n10960 ;
  assign n11088 = n11086 ^ x203 ;
  assign n11087 = n11086 ^ n11079 ;
  assign n11089 = n11088 ^ n11087 ;
  assign n11090 = n11084 & ~n11089 ;
  assign n11091 = n11090 ^ n11088 ;
  assign n11092 = n10964 ^ n9057 ;
  assign n11093 = n11092 ^ n10976 ;
  assign n11095 = n11093 ^ x202 ;
  assign n11094 = n11093 ^ n11086 ;
  assign n11096 = n11095 ^ n11094 ;
  assign n11097 = ~n11091 & n11096 ;
  assign n11098 = n11097 ^ n11095 ;
  assign n11100 = n11008 ^ x201 ;
  assign n11099 = n11093 ^ n11008 ;
  assign n11101 = n11100 ^ n11099 ;
  assign n11102 = n11098 & ~n11101 ;
  assign n11103 = n11102 ^ n11100 ;
  assign n11104 = ~n11009 & n11103 ;
  assign n11105 = n11104 ^ x200 ;
  assign n11005 = n11004 ^ n9111 ;
  assign n11006 = n11005 ^ n10995 ;
  assign n11106 = n11105 ^ n11006 ;
  assign n11120 = n11119 ^ n9870 ;
  assign n11121 = n11120 ^ x215 ;
  assign n11122 = n11121 ^ n11006 ;
  assign n11123 = n11122 ^ n11120 ;
  assign n11124 = ~n11106 & n11123 ;
  assign n11125 = n11124 ^ n11121 ;
  assign n11141 = n11140 ^ n11136 ;
  assign n11143 = n11141 ^ x214 ;
  assign n11142 = n11141 ^ n11120 ;
  assign n11144 = n11143 ^ n11142 ;
  assign n11145 = ~n11125 & n11144 ;
  assign n11146 = n11145 ^ n11143 ;
  assign n11150 = n11149 ^ n9245 ;
  assign n11162 = n11161 ^ n11150 ;
  assign n11164 = n11162 ^ x213 ;
  assign n11163 = n11162 ^ n11141 ;
  assign n11165 = n11164 ^ n11163 ;
  assign n11166 = ~n11146 & n11165 ;
  assign n11167 = n11166 ^ n11164 ;
  assign n11172 = n11171 ^ n9290 ;
  assign n11185 = n11184 ^ n11172 ;
  assign n11187 = n11185 ^ x212 ;
  assign n11186 = n11185 ^ n11162 ;
  assign n11188 = n11187 ^ n11186 ;
  assign n11189 = n11167 & ~n11188 ;
  assign n11190 = n11189 ^ n11187 ;
  assign n11195 = n11194 ^ n9335 ;
  assign n11208 = n11207 ^ n11195 ;
  assign n11210 = n11208 ^ x211 ;
  assign n11209 = n11208 ^ n11185 ;
  assign n11211 = n11210 ^ n11209 ;
  assign n11212 = n11190 & ~n11211 ;
  assign n11213 = n11212 ^ n11210 ;
  assign n11218 = n11217 ^ n9380 ;
  assign n11231 = n11230 ^ n11218 ;
  assign n11233 = n11231 ^ x210 ;
  assign n11232 = n11231 ^ n11208 ;
  assign n11234 = n11233 ^ n11232 ;
  assign n11235 = n11213 & ~n11234 ;
  assign n11236 = n11235 ^ n11233 ;
  assign n11250 = n11249 ^ n9425 ;
  assign n11251 = n11250 ^ n11245 ;
  assign n11253 = n11251 ^ x209 ;
  assign n11252 = n11251 ^ n11231 ;
  assign n11254 = n11253 ^ n11252 ;
  assign n11255 = ~n11236 & n11254 ;
  assign n11256 = n11255 ^ n11253 ;
  assign n11302 = n11251 ^ x208 ;
  assign n11303 = ~n11256 & n11302 ;
  assign n11304 = n11303 ^ x208 ;
  assign n11320 = n11319 ^ n11304 ;
  assign n11321 = n11319 ^ x223 ;
  assign n11322 = ~n11320 & n11321 ;
  assign n11323 = n11322 ^ x223 ;
  assign n11340 = n11339 ^ n11323 ;
  assign n11341 = n11337 ^ n11334 ;
  assign n11343 = n11330 ^ n11324 ;
  assign n11344 = ~n11329 & ~n11343 ;
  assign n11345 = n11344 ^ n11324 ;
  assign n11342 = n10748 ^ n10747 ;
  assign n11346 = n11345 ^ n11342 ;
  assign n11347 = n10092 & ~n11346 ;
  assign n11348 = n11347 ^ n10622 ;
  assign n11349 = n11348 ^ n9939 ;
  assign n11350 = n11349 ^ n11348 ;
  assign n11351 = n11350 ^ n11334 ;
  assign n11352 = ~n11341 & ~n11351 ;
  assign n11353 = n11352 ^ n11349 ;
  assign n11354 = n11353 ^ n9556 ;
  assign n11355 = n11354 ^ x222 ;
  assign n11356 = n11355 ^ n11354 ;
  assign n11357 = n11356 ^ n11323 ;
  assign n11358 = n11340 & n11357 ;
  assign n11359 = n11358 ^ n11355 ;
  assign n11369 = n10750 ^ n10749 ;
  assign n11365 = n10635 ^ n10622 ;
  assign n11364 = n11345 ^ n10635 ;
  assign n11366 = n11365 ^ n11364 ;
  assign n11367 = n11346 & ~n11366 ;
  assign n11368 = n11367 ^ n11365 ;
  assign n11370 = n11369 ^ n11368 ;
  assign n11371 = n11370 ^ n10635 ;
  assign n11372 = n10117 & n11371 ;
  assign n11373 = n11372 ^ n10635 ;
  assign n11360 = n11348 ^ n9556 ;
  assign n11361 = ~n11353 & n11360 ;
  assign n11362 = n11361 ^ n9556 ;
  assign n11363 = n11362 ^ n9599 ;
  assign n11374 = n11373 ^ n11363 ;
  assign n11376 = n11374 ^ x221 ;
  assign n11375 = n11374 ^ n11354 ;
  assign n11377 = n11376 ^ n11375 ;
  assign n11378 = n11359 & ~n11377 ;
  assign n11379 = n11378 ^ n11376 ;
  assign n11390 = n10752 ^ n10751 ;
  assign n11386 = n10660 ^ n10635 ;
  assign n11385 = n11369 ^ n10660 ;
  assign n11387 = n11386 ^ n11385 ;
  assign n11388 = ~n11368 & ~n11387 ;
  assign n11389 = n11388 ^ n11386 ;
  assign n11391 = n11390 ^ n11389 ;
  assign n11392 = n11391 ^ n10660 ;
  assign n11393 = ~n10138 & n11392 ;
  assign n11394 = n11393 ^ n10660 ;
  assign n11380 = n11373 ^ n11362 ;
  assign n11381 = n11373 ^ n9599 ;
  assign n11382 = n11380 & n11381 ;
  assign n11383 = n11382 ^ n9599 ;
  assign n11384 = n11383 ^ n9643 ;
  assign n11395 = n11394 ^ n11384 ;
  assign n11397 = n11395 ^ x220 ;
  assign n11396 = n11395 ^ n11374 ;
  assign n11398 = n11397 ^ n11396 ;
  assign n11399 = n11379 & ~n11398 ;
  assign n11400 = n11399 ^ n11397 ;
  assign n11412 = n11394 ^ n11383 ;
  assign n11413 = n11394 ^ n9643 ;
  assign n11414 = ~n11412 & ~n11413 ;
  assign n11415 = n11414 ^ n9643 ;
  assign n11416 = n11415 ^ n9676 ;
  assign n11407 = n10755 ^ n10753 ;
  assign n11401 = n10680 ^ n10158 ;
  assign n11403 = n11401 ^ n10660 ;
  assign n11402 = n11401 ^ n11390 ;
  assign n11404 = n11403 ^ n11402 ;
  assign n11405 = n11389 & n11404 ;
  assign n11406 = n11405 ^ n11403 ;
  assign n11408 = n11407 ^ n11406 ;
  assign n11409 = n11408 ^ n10680 ;
  assign n11410 = ~n10158 & ~n11409 ;
  assign n11411 = n11410 ^ n11408 ;
  assign n11417 = n11416 ^ n11411 ;
  assign n11419 = n11417 ^ x219 ;
  assign n11418 = n11417 ^ n11395 ;
  assign n11420 = n11419 ^ n11418 ;
  assign n11421 = n11400 & ~n11420 ;
  assign n11422 = n11421 ^ n11419 ;
  assign n11430 = n11407 ^ n11401 ;
  assign n11431 = ~n11406 & n11430 ;
  assign n11429 = n11401 ^ n10700 ;
  assign n11432 = n11431 ^ n11429 ;
  assign n11428 = n10757 ^ n10756 ;
  assign n11433 = n11432 ^ n11428 ;
  assign n11434 = n11433 ^ n10700 ;
  assign n11435 = n10179 & ~n11434 ;
  assign n11436 = n11435 ^ n10700 ;
  assign n11423 = n11415 ^ n11411 ;
  assign n11424 = n11411 ^ n9676 ;
  assign n11425 = n11423 & n11424 ;
  assign n11426 = n11425 ^ n9676 ;
  assign n11427 = n11426 ^ n9730 ;
  assign n11437 = n11436 ^ n11427 ;
  assign n11439 = n11437 ^ x218 ;
  assign n11438 = n11437 ^ n11417 ;
  assign n11440 = n11439 ^ n11438 ;
  assign n11441 = n11422 & ~n11440 ;
  assign n11442 = n11441 ^ n11439 ;
  assign n11257 = n11256 ^ x208 ;
  assign n11258 = n11103 ^ x200 ;
  assign n11268 = ~n11266 & ~n11267 ;
  assign n11269 = n11077 ^ x204 ;
  assign n11270 = n11268 & n11269 ;
  assign n11271 = n11084 ^ x203 ;
  assign n11272 = ~n11270 & n11271 ;
  assign n11273 = n11091 ^ x202 ;
  assign n11274 = n11272 & ~n11273 ;
  assign n11275 = n11098 ^ x201 ;
  assign n11276 = ~n11274 & ~n11275 ;
  assign n11277 = n11258 & ~n11276 ;
  assign n11278 = n11105 ^ x215 ;
  assign n11279 = n11278 ^ n11006 ;
  assign n11280 = ~n11277 & n11279 ;
  assign n11281 = n11125 ^ x214 ;
  assign n11282 = n11280 & n11281 ;
  assign n11283 = n11146 ^ x213 ;
  assign n11284 = n11282 & n11283 ;
  assign n11285 = n11167 ^ x212 ;
  assign n11286 = n11284 & ~n11285 ;
  assign n11287 = n11190 ^ x211 ;
  assign n11288 = n11286 & ~n11287 ;
  assign n11289 = n11213 ^ x210 ;
  assign n11290 = n11288 & ~n11289 ;
  assign n11291 = n11236 ^ x209 ;
  assign n11292 = ~n11290 & ~n11291 ;
  assign n11444 = n11257 & ~n11292 ;
  assign n11445 = n11304 ^ x223 ;
  assign n11446 = n11445 ^ n11319 ;
  assign n11447 = n11444 & n11446 ;
  assign n11448 = n11340 ^ x222 ;
  assign n11449 = n11447 & ~n11448 ;
  assign n11450 = n11359 ^ x221 ;
  assign n11451 = n11449 & ~n11450 ;
  assign n11452 = n11379 ^ x220 ;
  assign n11453 = n11451 & ~n11452 ;
  assign n11454 = n11400 ^ x219 ;
  assign n11455 = n11453 & ~n11454 ;
  assign n11456 = n11422 ^ x218 ;
  assign n11457 = n11455 & ~n11456 ;
  assign n11519 = n11457 ^ n11437 ;
  assign n11520 = n11442 & n11519 ;
  assign n11517 = n11457 ^ n11442 ;
  assign n11518 = x217 & n11517 ;
  assign n11521 = n11520 ^ n11518 ;
  assign n11513 = n9730 ^ x216 ;
  assign n11512 = n10785 ^ n9807 ;
  assign n11514 = n11513 ^ n11512 ;
  assign n11507 = n11428 ^ n10700 ;
  assign n11508 = n11432 & n11507 ;
  assign n11505 = n10760 ^ n10758 ;
  assign n11504 = n11428 ^ n10785 ;
  assign n11506 = n11505 ^ n11504 ;
  assign n11509 = n11508 ^ n11506 ;
  assign n11510 = n11509 ^ n10785 ;
  assign n11511 = ~n10229 & ~n11510 ;
  assign n11515 = n11514 ^ n11511 ;
  assign n11501 = n11436 ^ n11426 ;
  assign n11502 = n11436 ^ n9730 ;
  assign n11503 = ~n11501 & ~n11502 ;
  assign n11516 = n11515 ^ n11503 ;
  assign n11522 = n11521 ^ n11516 ;
  assign n11443 = n11442 ^ x217 ;
  assign n11458 = n11457 ^ n11443 ;
  assign n11459 = n11458 ^ n10885 ;
  assign n11461 = n10823 ^ n9897 ;
  assign n11460 = n11456 ^ n11455 ;
  assign n11462 = n11461 ^ n11460 ;
  assign n11463 = n11454 ^ n11453 ;
  assign n11464 = n11463 ^ n10840 ;
  assign n11466 = n11452 ^ n11451 ;
  assign n11465 = n10815 ^ n10789 ;
  assign n11467 = n11466 ^ n11465 ;
  assign n11469 = n10811 ^ n10794 ;
  assign n11470 = n11469 ^ n10792 ;
  assign n11468 = n11450 ^ n11449 ;
  assign n11471 = n11470 ^ n11468 ;
  assign n11473 = n11448 ^ n11447 ;
  assign n11472 = n10809 ^ n10798 ;
  assign n11474 = n11473 ^ n11472 ;
  assign n11477 = n10805 ^ n10804 ;
  assign n11293 = n11292 ^ n11257 ;
  assign n11475 = n10800 ^ n9533 ;
  assign n11476 = ~n11293 & n11475 ;
  assign n11478 = n11477 ^ n11476 ;
  assign n11479 = n11446 ^ n11444 ;
  assign n11480 = n11479 ^ n11476 ;
  assign n11481 = n11478 & ~n11480 ;
  assign n11482 = n11481 ^ n11477 ;
  assign n11483 = n11482 ^ n11472 ;
  assign n11484 = ~n11474 & ~n11483 ;
  assign n11485 = n11484 ^ n11473 ;
  assign n11486 = n11485 ^ n11468 ;
  assign n11487 = ~n11471 & ~n11486 ;
  assign n11488 = n11487 ^ n11470 ;
  assign n11489 = n11488 ^ n11465 ;
  assign n11490 = ~n11467 & ~n11489 ;
  assign n11491 = n11490 ^ n11466 ;
  assign n11492 = n11491 ^ n11463 ;
  assign n11493 = n11464 & ~n11492 ;
  assign n11494 = n11493 ^ n10840 ;
  assign n11495 = n11494 ^ n11460 ;
  assign n11496 = ~n11462 & ~n11495 ;
  assign n11497 = n11496 ^ n11461 ;
  assign n11498 = n11497 ^ n11458 ;
  assign n11499 = n11459 & ~n11498 ;
  assign n11500 = n11499 ^ n10885 ;
  assign n11523 = n11522 ^ n11500 ;
  assign n11524 = n11298 ^ n10892 ;
  assign n11525 = n11524 ^ n11298 ;
  assign n11526 = n11525 ^ n11500 ;
  assign n11527 = n11523 & ~n11526 ;
  assign n11528 = n11527 ^ n11524 ;
  assign n11529 = n11301 & ~n11528 ;
  assign n11299 = n11298 ^ n10910 ;
  assign n11530 = n11529 ^ n11299 ;
  assign n11531 = n11016 ^ x198 ;
  assign n11532 = n11531 ^ n11014 ;
  assign n11533 = n11532 ^ n10910 ;
  assign n11534 = n11530 & n11533 ;
  assign n11536 = n11535 ^ n11534 ;
  assign n11539 = n11023 ^ x197 ;
  assign n11537 = n10941 ^ n10925 ;
  assign n11538 = n11537 ^ n10941 ;
  assign n11540 = n11539 ^ n11538 ;
  assign n11541 = ~n11536 & ~n11540 ;
  assign n11542 = n11541 ^ n11537 ;
  assign n11545 = n10957 ^ n10941 ;
  assign n11543 = n11029 ^ x196 ;
  assign n11544 = n11543 ^ n10957 ;
  assign n11546 = n11545 ^ n11544 ;
  assign n11547 = n11542 & n11546 ;
  assign n11548 = n11547 ^ n11545 ;
  assign n11551 = n10973 ^ n10957 ;
  assign n11549 = n11035 ^ x195 ;
  assign n11550 = n11549 ^ n10973 ;
  assign n11552 = n11551 ^ n11550 ;
  assign n11553 = ~n11548 & ~n11552 ;
  assign n11554 = n11553 ^ n11551 ;
  assign n11555 = n11041 ^ x194 ;
  assign n11563 = n11555 ^ n10973 ;
  assign n11564 = ~n11554 & ~n11563 ;
  assign n11565 = n11564 ^ n10973 ;
  assign n11566 = n11565 ^ n11259 ;
  assign n11567 = ~n11562 & n11566 ;
  assign n11561 = n11558 ^ n10988 ;
  assign n11568 = n11567 ^ n11561 ;
  assign n11569 = n11560 & n11568 ;
  assign n11570 = n11569 ^ n11559 ;
  assign n11572 = n11571 ^ n11570 ;
  assign n11573 = n11127 ^ n11112 ;
  assign n11576 = n11573 ^ n11570 ;
  assign n11577 = n11572 & ~n11576 ;
  assign n11574 = n11573 ^ n11133 ;
  assign n11578 = n11577 ^ n11574 ;
  assign n11581 = n11158 ^ n11133 ;
  assign n11579 = n11265 ^ n11264 ;
  assign n11580 = n11579 ^ n11158 ;
  assign n11582 = n11581 ^ n11580 ;
  assign n11583 = ~n11578 & n11582 ;
  assign n11584 = n11583 ^ n11581 ;
  assign n11619 = n11585 ^ n11584 ;
  assign n11948 = n11279 ^ n11277 ;
  assign n11775 = n11311 ^ n10324 ;
  assign n11776 = n11775 ^ n11242 ;
  assign n11587 = n11181 ^ n11158 ;
  assign n11586 = n11585 ^ n11181 ;
  assign n11588 = n11587 ^ n11586 ;
  assign n11589 = n11584 & n11588 ;
  assign n11590 = n11589 ^ n11587 ;
  assign n11593 = n11204 ^ n11181 ;
  assign n11591 = n11269 ^ n11268 ;
  assign n11592 = n11591 ^ n11204 ;
  assign n11594 = n11593 ^ n11592 ;
  assign n11595 = ~n11590 & ~n11594 ;
  assign n11596 = n11595 ^ n11593 ;
  assign n11599 = n11227 ^ n11204 ;
  assign n11597 = n11271 ^ n11270 ;
  assign n11598 = n11597 ^ n11227 ;
  assign n11600 = n11599 ^ n11598 ;
  assign n11601 = ~n11596 & n11600 ;
  assign n11602 = n11601 ^ n11599 ;
  assign n11763 = n11242 ^ n11227 ;
  assign n11603 = n11273 ^ n11272 ;
  assign n11762 = n11603 ^ n11242 ;
  assign n11764 = n11763 ^ n11762 ;
  assign n11765 = ~n11602 & ~n11764 ;
  assign n11766 = n11765 ^ n11763 ;
  assign n11767 = n11275 ^ n11274 ;
  assign n11773 = n11767 ^ n11242 ;
  assign n11774 = ~n11766 & n11773 ;
  assign n11777 = n11776 ^ n11774 ;
  assign n11778 = n11276 ^ n11258 ;
  assign n11945 = n11778 ^ n11775 ;
  assign n11946 = n11777 & ~n11945 ;
  assign n11947 = n11946 ^ n11778 ;
  assign n11949 = n11948 ^ n11947 ;
  assign n12664 = n11949 ^ n11331 ;
  assign n11768 = n11767 ^ n11766 ;
  assign n11604 = n11603 ^ n11602 ;
  assign n12418 = n11768 ^ n11604 ;
  assign n11294 = n9533 & n11293 ;
  assign n11295 = n11294 ^ n10800 ;
  assign n11296 = n11295 ^ n9091 ;
  assign n11803 = x359 & ~n11296 ;
  assign n11672 = ~n9091 & n11295 ;
  assign n11674 = n11672 ^ n9128 ;
  assign n11670 = n10803 & n11480 ;
  assign n11671 = n11670 ^ n11477 ;
  assign n11802 = n11674 ^ n11671 ;
  assign n11804 = n11803 ^ n11802 ;
  assign n11673 = n11672 ^ n11671 ;
  assign n11675 = ~n11673 & n11674 ;
  assign n11676 = n11675 ^ n9128 ;
  assign n11678 = n11676 ^ n9166 ;
  assign n11667 = n11482 ^ n11473 ;
  assign n11668 = n10797 & ~n11667 ;
  assign n11669 = n11668 ^ n11472 ;
  assign n11805 = n11678 ^ n11669 ;
  assign n11806 = n11805 ^ x358 ;
  assign n11807 = n11806 ^ n11803 ;
  assign n11808 = n11807 ^ n11805 ;
  assign n11809 = ~n11804 & n11808 ;
  assign n11810 = n11809 ^ n11806 ;
  assign n11677 = n11676 ^ n11669 ;
  assign n11679 = ~n11677 & n11678 ;
  assign n11680 = n11679 ^ n9166 ;
  assign n11682 = n11680 ^ n9212 ;
  assign n11665 = n10794 & n11486 ;
  assign n11666 = n11665 ^ n11470 ;
  assign n11811 = n11682 ^ n11666 ;
  assign n11813 = n11811 ^ x357 ;
  assign n11812 = n11811 ^ n11805 ;
  assign n11814 = n11813 ^ n11812 ;
  assign n11815 = ~n11810 & n11814 ;
  assign n11816 = n11815 ^ n11813 ;
  assign n11681 = n11680 ^ n11666 ;
  assign n11683 = ~n11681 & ~n11682 ;
  assign n11684 = n11683 ^ n9212 ;
  assign n11686 = n11684 ^ n9256 ;
  assign n11662 = n11488 ^ n11466 ;
  assign n11663 = ~n9938 & ~n11662 ;
  assign n11664 = n11663 ^ n11465 ;
  assign n11817 = n11686 ^ n11664 ;
  assign n11819 = n11817 ^ x356 ;
  assign n11818 = n11817 ^ n11811 ;
  assign n11820 = n11819 ^ n11818 ;
  assign n11821 = n11816 & ~n11820 ;
  assign n11822 = n11821 ^ n11819 ;
  assign n12023 = n11822 ^ x355 ;
  assign n12017 = n11810 ^ x357 ;
  assign n11297 = n11296 ^ x359 ;
  assign n12018 = n11804 ^ x358 ;
  assign n12019 = ~n11297 & n12018 ;
  assign n12020 = n12017 & n12019 ;
  assign n12021 = n11816 ^ x356 ;
  assign n12022 = n12020 & ~n12021 ;
  assign n12225 = n12023 ^ n12022 ;
  assign n11624 = n11579 ^ n11578 ;
  assign n12226 = n12225 ^ n11624 ;
  assign n12228 = n12021 ^ n12020 ;
  assign n12250 = n12228 ^ n11624 ;
  assign n12227 = n11573 ^ n11572 ;
  assign n12229 = n12228 ^ n12227 ;
  assign n12240 = n12019 ^ n12017 ;
  assign n12231 = n11565 ^ n11562 ;
  assign n12241 = n12240 ^ n12231 ;
  assign n12230 = n12018 ^ n11297 ;
  assign n12232 = n12231 ^ n12230 ;
  assign n11950 = n11324 & ~n11949 ;
  assign n11951 = n11950 ^ n11331 ;
  assign n11769 = n11768 ^ n11242 ;
  assign n11770 = n10450 & ~n11769 ;
  assign n11771 = n11770 ^ n11242 ;
  assign n11605 = n11604 ^ n11227 ;
  assign n11606 = ~n11220 & n11605 ;
  assign n11607 = n11606 ^ n11227 ;
  assign n11608 = n11607 ^ n10014 ;
  assign n11609 = n11597 ^ n11596 ;
  assign n11610 = n11609 ^ n11204 ;
  assign n11611 = n11197 & ~n11610 ;
  assign n11612 = n11611 ^ n11204 ;
  assign n11613 = n11612 ^ n9994 ;
  assign n11614 = n11591 ^ n11590 ;
  assign n11615 = n11614 ^ n11181 ;
  assign n11616 = n11174 & n11615 ;
  assign n11617 = n11616 ^ n11181 ;
  assign n11618 = n11617 ^ n9973 ;
  assign n11620 = n11619 ^ n11158 ;
  assign n11621 = ~n11151 & n11620 ;
  assign n11622 = n11621 ^ n11158 ;
  assign n11623 = n11622 ^ n9952 ;
  assign n11625 = n11624 ^ n11133 ;
  assign n11626 = n11130 & ~n11625 ;
  assign n11627 = n11626 ^ n11133 ;
  assign n11628 = n11627 ^ n9875 ;
  assign n11727 = ~n10981 & ~n11566 ;
  assign n11728 = n11727 ^ n10988 ;
  assign n11556 = n11555 ^ n11554 ;
  assign n11629 = n11556 ^ n10973 ;
  assign n11630 = n10966 & n11629 ;
  assign n11631 = n11630 ^ n10973 ;
  assign n11632 = n11631 ^ n9693 ;
  assign n11633 = n11549 ^ n11548 ;
  assign n11634 = n11633 ^ n10957 ;
  assign n11635 = n10950 & n11634 ;
  assign n11636 = n11635 ^ n10957 ;
  assign n11637 = n11636 ^ n9654 ;
  assign n11638 = n11543 ^ n11542 ;
  assign n11639 = n11638 ^ n10941 ;
  assign n11640 = ~n10934 & n11639 ;
  assign n11641 = n11640 ^ n10941 ;
  assign n11642 = n11641 ^ n9610 ;
  assign n11643 = n11539 ^ n11536 ;
  assign n11644 = n11643 ^ n10925 ;
  assign n11645 = n10918 & n11644 ;
  assign n11646 = n11645 ^ n10925 ;
  assign n11647 = n11646 ^ n9567 ;
  assign n11648 = n11532 ^ n11530 ;
  assign n11649 = n11648 ^ n10910 ;
  assign n11650 = n10907 & n11649 ;
  assign n11651 = n11650 ^ n10910 ;
  assign n11652 = n11651 ^ n9522 ;
  assign n11653 = ~n9886 & ~n11523 ;
  assign n11654 = n11653 ^ n10892 ;
  assign n11655 = n11654 ^ n9436 ;
  assign n11685 = n11684 ^ n11664 ;
  assign n11687 = n11685 & ~n11686 ;
  assign n11688 = n11687 ^ n9256 ;
  assign n11660 = n9934 & n11492 ;
  assign n11661 = n11660 ^ n10840 ;
  assign n11689 = n11688 ^ n11661 ;
  assign n11690 = n11688 ^ n9301 ;
  assign n11691 = n11689 & n11690 ;
  assign n11692 = n11691 ^ n9301 ;
  assign n11658 = n10822 & n11495 ;
  assign n11659 = n11658 ^ n11461 ;
  assign n11693 = n11692 ^ n11659 ;
  assign n11694 = n11692 ^ n9346 ;
  assign n11695 = ~n11693 & ~n11694 ;
  assign n11696 = n11695 ^ n9346 ;
  assign n11656 = n9930 & n11498 ;
  assign n11657 = n11656 ^ n10885 ;
  assign n11697 = n11696 ^ n11657 ;
  assign n11698 = n11696 ^ n9391 ;
  assign n11699 = n11697 & n11698 ;
  assign n11700 = n11699 ^ n9391 ;
  assign n11701 = n11700 ^ n11654 ;
  assign n11702 = n11655 & ~n11701 ;
  assign n11703 = n11702 ^ n9436 ;
  assign n11704 = n11703 ^ n9480 ;
  assign n11705 = n11528 ^ n11300 ;
  assign n11706 = n11705 ^ n10834 ;
  assign n11707 = n10837 & ~n11706 ;
  assign n11708 = n11707 ^ n10834 ;
  assign n11709 = n11708 ^ n11703 ;
  assign n11710 = n11704 & n11709 ;
  assign n11711 = n11710 ^ n9480 ;
  assign n11712 = n11711 ^ n11651 ;
  assign n11713 = ~n11652 & n11712 ;
  assign n11714 = n11713 ^ n9522 ;
  assign n11715 = n11714 ^ n11646 ;
  assign n11716 = ~n11647 & ~n11715 ;
  assign n11717 = n11716 ^ n9567 ;
  assign n11718 = n11717 ^ n11641 ;
  assign n11719 = n11642 & n11718 ;
  assign n11720 = n11719 ^ n9610 ;
  assign n11721 = n11720 ^ n11636 ;
  assign n11722 = ~n11637 & n11721 ;
  assign n11723 = n11722 ^ n9654 ;
  assign n11724 = n11723 ^ n11631 ;
  assign n11725 = n11632 & ~n11724 ;
  assign n11726 = n11725 ^ n9693 ;
  assign n11729 = n11728 ^ n11726 ;
  assign n11730 = ~n11003 & ~n11568 ;
  assign n11731 = n11730 ^ n11559 ;
  assign n11732 = n11731 ^ n9741 ;
  assign n11733 = n11732 ^ n11726 ;
  assign n11734 = n11733 ^ n11731 ;
  assign n11735 = ~n11729 & n11734 ;
  assign n11736 = n11735 ^ n11732 ;
  assign n11737 = ~n11127 & n11572 ;
  assign n11738 = n11737 ^ n11112 ;
  assign n11740 = n11738 ^ n9822 ;
  assign n11739 = n11738 ^ n11731 ;
  assign n11741 = n11740 ^ n11739 ;
  assign n11742 = n11736 & ~n11741 ;
  assign n11743 = n11742 ^ n11740 ;
  assign n11744 = n11738 ^ n10241 ;
  assign n11745 = n11743 & n11744 ;
  assign n11746 = n11745 ^ n10241 ;
  assign n11747 = n11746 ^ n11627 ;
  assign n11748 = ~n11628 & ~n11747 ;
  assign n11749 = n11748 ^ n9875 ;
  assign n11750 = n11749 ^ n11622 ;
  assign n11751 = ~n11623 & n11750 ;
  assign n11752 = n11751 ^ n9952 ;
  assign n11753 = n11752 ^ n11617 ;
  assign n11754 = n11618 & ~n11753 ;
  assign n11755 = n11754 ^ n9973 ;
  assign n11756 = n11755 ^ n11612 ;
  assign n11757 = ~n11613 & n11756 ;
  assign n11758 = n11757 ^ n9994 ;
  assign n11759 = n11758 ^ n11607 ;
  assign n11760 = n11608 & ~n11759 ;
  assign n11761 = n11760 ^ n10014 ;
  assign n11772 = n11771 ^ n11761 ;
  assign n11779 = n11778 ^ n11777 ;
  assign n11780 = n11779 ^ n11311 ;
  assign n11781 = n10324 & ~n11780 ;
  assign n11782 = n11781 ^ n11779 ;
  assign n11783 = n11782 ^ n10035 ;
  assign n11784 = n11783 ^ n11761 ;
  assign n11785 = n11784 ^ n11782 ;
  assign n11786 = n11772 & ~n11785 ;
  assign n11787 = n11786 ^ n11783 ;
  assign n11941 = n11782 ^ n10050 ;
  assign n11942 = n11787 & n11941 ;
  assign n11943 = n11942 ^ n10050 ;
  assign n11944 = n11943 ^ n10616 ;
  assign n11952 = n11951 ^ n11944 ;
  assign n11788 = n11787 ^ n10050 ;
  assign n11789 = n11788 ^ x383 ;
  assign n11790 = n11761 ^ n10035 ;
  assign n11791 = n11790 ^ n11771 ;
  assign n11792 = n11791 ^ x368 ;
  assign n11921 = n11755 ^ n9994 ;
  assign n11922 = n11921 ^ n11612 ;
  assign n11793 = n11752 ^ n9973 ;
  assign n11794 = n11793 ^ n11617 ;
  assign n11795 = n11794 ^ x371 ;
  assign n11892 = n11736 ^ n9822 ;
  assign n11796 = n11726 ^ n9741 ;
  assign n11797 = n11796 ^ n11728 ;
  assign n11798 = n11797 ^ x360 ;
  assign n11882 = n11723 ^ n9693 ;
  assign n11883 = n11882 ^ n11631 ;
  assign n11799 = n11720 ^ n9654 ;
  assign n11800 = n11799 ^ n11636 ;
  assign n11801 = n11800 ^ x362 ;
  assign n11823 = n11690 ^ n11661 ;
  assign n11825 = n11823 ^ x355 ;
  assign n11824 = n11823 ^ n11817 ;
  assign n11826 = n11825 ^ n11824 ;
  assign n11827 = n11822 & ~n11826 ;
  assign n11828 = n11827 ^ n11825 ;
  assign n11829 = n11694 ^ n11659 ;
  assign n11831 = n11829 ^ x354 ;
  assign n11830 = n11829 ^ n11823 ;
  assign n11832 = n11831 ^ n11830 ;
  assign n11833 = n11828 & ~n11832 ;
  assign n11834 = n11833 ^ n11831 ;
  assign n11835 = n11698 ^ n11657 ;
  assign n11837 = n11835 ^ x353 ;
  assign n11836 = n11835 ^ n11829 ;
  assign n11838 = n11837 ^ n11836 ;
  assign n11839 = n11834 & ~n11838 ;
  assign n11840 = n11839 ^ n11837 ;
  assign n11841 = n11700 ^ n9436 ;
  assign n11842 = n11841 ^ n11654 ;
  assign n11844 = n11842 ^ x352 ;
  assign n11843 = n11842 ^ n11835 ;
  assign n11845 = n11844 ^ n11843 ;
  assign n11846 = ~n11840 & n11845 ;
  assign n11847 = n11846 ^ n11844 ;
  assign n11848 = n11708 ^ n11704 ;
  assign n11850 = n11848 ^ x367 ;
  assign n11849 = n11848 ^ n11842 ;
  assign n11851 = n11850 ^ n11849 ;
  assign n11852 = n11847 & ~n11851 ;
  assign n11853 = n11852 ^ n11850 ;
  assign n11854 = n11711 ^ n9522 ;
  assign n11855 = n11854 ^ n11651 ;
  assign n11857 = n11855 ^ x366 ;
  assign n11856 = n11855 ^ n11848 ;
  assign n11858 = n11857 ^ n11856 ;
  assign n11859 = ~n11853 & n11858 ;
  assign n11860 = n11859 ^ n11857 ;
  assign n11861 = n11714 ^ n9567 ;
  assign n11862 = n11861 ^ n11646 ;
  assign n11864 = n11862 ^ x365 ;
  assign n11863 = n11862 ^ n11855 ;
  assign n11865 = n11864 ^ n11863 ;
  assign n11866 = ~n11860 & n11865 ;
  assign n11867 = n11866 ^ n11864 ;
  assign n11868 = n11717 ^ n9610 ;
  assign n11869 = n11868 ^ n11641 ;
  assign n11871 = n11869 ^ x364 ;
  assign n11870 = n11869 ^ n11862 ;
  assign n11872 = n11871 ^ n11870 ;
  assign n11873 = ~n11867 & n11872 ;
  assign n11874 = n11873 ^ n11871 ;
  assign n11876 = n11800 ^ x363 ;
  assign n11875 = n11869 ^ n11800 ;
  assign n11877 = n11876 ^ n11875 ;
  assign n11878 = ~n11874 & n11877 ;
  assign n11879 = n11878 ^ n11876 ;
  assign n11880 = n11801 & ~n11879 ;
  assign n11881 = n11880 ^ x362 ;
  assign n11884 = n11883 ^ n11881 ;
  assign n11886 = n11797 ^ x361 ;
  assign n11885 = n11881 ^ n11797 ;
  assign n11887 = n11886 ^ n11885 ;
  assign n11888 = n11884 & n11887 ;
  assign n11889 = n11888 ^ n11886 ;
  assign n11890 = ~n11798 & n11889 ;
  assign n11891 = n11890 ^ x360 ;
  assign n11893 = n11892 ^ n11891 ;
  assign n11894 = n11743 ^ n10241 ;
  assign n11895 = n11894 ^ x375 ;
  assign n11896 = n11895 ^ n11891 ;
  assign n11897 = n11896 ^ n11894 ;
  assign n11898 = ~n11893 & n11897 ;
  assign n11899 = n11898 ^ n11895 ;
  assign n11900 = n11746 ^ n9875 ;
  assign n11901 = n11900 ^ n11627 ;
  assign n11903 = n11901 ^ x374 ;
  assign n11902 = n11901 ^ n11894 ;
  assign n11904 = n11903 ^ n11902 ;
  assign n11905 = n11899 & ~n11904 ;
  assign n11906 = n11905 ^ n11903 ;
  assign n11907 = n11749 ^ n9952 ;
  assign n11908 = n11907 ^ n11622 ;
  assign n11910 = n11908 ^ x373 ;
  assign n11909 = n11908 ^ n11901 ;
  assign n11911 = n11910 ^ n11909 ;
  assign n11912 = n11906 & ~n11911 ;
  assign n11913 = n11912 ^ n11910 ;
  assign n11915 = n11794 ^ x372 ;
  assign n11914 = n11908 ^ n11794 ;
  assign n11916 = n11915 ^ n11914 ;
  assign n11917 = ~n11913 & n11916 ;
  assign n11918 = n11917 ^ n11915 ;
  assign n11919 = ~n11795 & n11918 ;
  assign n11920 = n11919 ^ x371 ;
  assign n11923 = n11922 ^ n11920 ;
  assign n11924 = n11758 ^ n10014 ;
  assign n11925 = n11924 ^ n11607 ;
  assign n11926 = n11925 ^ x370 ;
  assign n11927 = n11926 ^ n11920 ;
  assign n11928 = n11927 ^ n11925 ;
  assign n11929 = ~n11923 & n11928 ;
  assign n11930 = n11929 ^ n11926 ;
  assign n11932 = n11791 ^ x369 ;
  assign n11931 = n11925 ^ n11791 ;
  assign n11933 = n11932 ^ n11931 ;
  assign n11934 = n11930 & ~n11933 ;
  assign n11935 = n11934 ^ n11932 ;
  assign n11936 = ~n11792 & n11935 ;
  assign n11937 = n11936 ^ x368 ;
  assign n11938 = n11937 ^ n11788 ;
  assign n11939 = n11789 & ~n11938 ;
  assign n11940 = n11939 ^ x383 ;
  assign n11953 = n11952 ^ n11940 ;
  assign n11965 = n11281 ^ n11280 ;
  assign n11959 = n11346 ^ n10622 ;
  assign n11960 = n11959 ^ n11331 ;
  assign n11961 = n11960 ^ n11959 ;
  assign n11962 = n11961 ^ n11947 ;
  assign n11963 = n11949 & n11962 ;
  assign n11964 = n11963 ^ n11960 ;
  assign n11966 = n11965 ^ n11964 ;
  assign n11967 = n11966 ^ n11346 ;
  assign n11968 = ~n10622 & ~n11967 ;
  assign n11969 = n11968 ^ n11346 ;
  assign n11954 = n11951 ^ n11943 ;
  assign n11955 = n11951 ^ n10616 ;
  assign n11956 = n11954 & n11955 ;
  assign n11957 = n11956 ^ n10616 ;
  assign n11958 = n11957 ^ n10092 ;
  assign n11970 = n11969 ^ n11958 ;
  assign n11971 = n11970 ^ x382 ;
  assign n11972 = n11971 ^ n11940 ;
  assign n11973 = n11972 ^ n11970 ;
  assign n11974 = n11953 & n11973 ;
  assign n11975 = n11974 ^ n11971 ;
  assign n11981 = n11283 ^ n11282 ;
  assign n11983 = n11981 ^ n11959 ;
  assign n11982 = n11981 ^ n11965 ;
  assign n11984 = n11983 ^ n11982 ;
  assign n11985 = n11964 & n11984 ;
  assign n11986 = n11985 ^ n11983 ;
  assign n11987 = n10635 & n11986 ;
  assign n11988 = n11987 ^ n11370 ;
  assign n11976 = n11969 ^ n11957 ;
  assign n11977 = n11969 ^ n10092 ;
  assign n11978 = n11976 & ~n11977 ;
  assign n11979 = n11978 ^ n10092 ;
  assign n11980 = n11979 ^ n10117 ;
  assign n11989 = n11988 ^ n11980 ;
  assign n11991 = n11989 ^ x381 ;
  assign n11990 = n11989 ^ n11970 ;
  assign n11992 = n11991 ^ n11990 ;
  assign n11993 = n11975 & ~n11992 ;
  assign n11994 = n11993 ^ n11991 ;
  assign n12005 = n11285 ^ n11284 ;
  assign n12001 = n11391 ^ n11370 ;
  assign n12000 = n11981 ^ n11391 ;
  assign n12002 = n12001 ^ n12000 ;
  assign n12003 = ~n11986 & n12002 ;
  assign n12004 = n12003 ^ n12001 ;
  assign n12006 = n12005 ^ n12004 ;
  assign n12007 = n12006 ^ n11391 ;
  assign n12008 = n10660 & ~n12007 ;
  assign n12009 = n12008 ^ n11391 ;
  assign n11995 = n11988 ^ n11979 ;
  assign n11996 = n11988 ^ n10117 ;
  assign n11997 = ~n11995 & n11996 ;
  assign n11998 = n11997 ^ n10117 ;
  assign n11999 = n11998 ^ n10138 ;
  assign n12010 = n12009 ^ n11999 ;
  assign n12012 = n12010 ^ x380 ;
  assign n12011 = n12010 ^ n11989 ;
  assign n12013 = n12012 ^ n12011 ;
  assign n12014 = ~n11994 & n12013 ;
  assign n12015 = n12014 ^ n12012 ;
  assign n12016 = n12015 ^ x379 ;
  assign n12024 = ~n12022 & n12023 ;
  assign n12025 = n11828 ^ x354 ;
  assign n12026 = ~n12024 & ~n12025 ;
  assign n12027 = n11834 ^ x353 ;
  assign n12028 = ~n12026 & n12027 ;
  assign n12029 = n11840 ^ x352 ;
  assign n12030 = ~n12028 & n12029 ;
  assign n12031 = n11847 ^ x367 ;
  assign n12032 = n12030 & ~n12031 ;
  assign n12033 = n11853 ^ x366 ;
  assign n12034 = ~n12032 & ~n12033 ;
  assign n12035 = n11860 ^ x365 ;
  assign n12036 = ~n12034 & n12035 ;
  assign n12037 = n11867 ^ x364 ;
  assign n12038 = ~n12036 & ~n12037 ;
  assign n12039 = n11874 ^ x363 ;
  assign n12040 = n12038 & ~n12039 ;
  assign n12041 = n11879 ^ x362 ;
  assign n12042 = ~n12040 & n12041 ;
  assign n12043 = n11884 ^ x361 ;
  assign n12044 = ~n12042 & n12043 ;
  assign n12045 = n11889 ^ x360 ;
  assign n12046 = ~n12044 & ~n12045 ;
  assign n12047 = n11891 ^ x375 ;
  assign n12048 = n12047 ^ n11892 ;
  assign n12049 = n12046 & n12048 ;
  assign n12050 = n11899 ^ x374 ;
  assign n12051 = ~n12049 & n12050 ;
  assign n12052 = n11906 ^ x373 ;
  assign n12053 = n12051 & n12052 ;
  assign n12054 = n11913 ^ x372 ;
  assign n12055 = n12053 & ~n12054 ;
  assign n12056 = n11918 ^ x371 ;
  assign n12057 = n12055 & n12056 ;
  assign n12058 = n11923 ^ x370 ;
  assign n12059 = ~n12057 & n12058 ;
  assign n12060 = n11930 ^ x369 ;
  assign n12061 = ~n12059 & n12060 ;
  assign n12062 = n11935 ^ x368 ;
  assign n12063 = ~n12061 & ~n12062 ;
  assign n12064 = n11937 ^ x383 ;
  assign n12065 = n12064 ^ n11788 ;
  assign n12066 = n12063 & n12065 ;
  assign n12067 = n11953 ^ x382 ;
  assign n12068 = ~n12066 & n12067 ;
  assign n12069 = n11975 ^ x381 ;
  assign n12070 = n12068 & n12069 ;
  assign n12071 = n11994 ^ x380 ;
  assign n12072 = ~n12070 & n12071 ;
  assign n12073 = ~n12016 & n12072 ;
  assign n12079 = n11287 ^ n11286 ;
  assign n12081 = n12079 ^ n11391 ;
  assign n12080 = n12079 ^ n12005 ;
  assign n12082 = n12081 ^ n12080 ;
  assign n12083 = n12004 & ~n12082 ;
  assign n12084 = n12083 ^ n12081 ;
  assign n12085 = ~n11401 & ~n12084 ;
  assign n12086 = n12085 ^ n11408 ;
  assign n12074 = n12009 ^ n11998 ;
  assign n12075 = n12009 ^ n10138 ;
  assign n12076 = ~n12074 & ~n12075 ;
  assign n12077 = n12076 ^ n10138 ;
  assign n12078 = n12077 ^ n10158 ;
  assign n12087 = n12086 ^ n12078 ;
  assign n12089 = n12087 ^ x379 ;
  assign n12088 = n12087 ^ n12010 ;
  assign n12090 = n12089 ^ n12088 ;
  assign n12091 = n12015 & ~n12090 ;
  assign n12092 = n12091 ^ n12089 ;
  assign n12093 = n12092 ^ x378 ;
  assign n12187 = ~n12073 & n12093 ;
  assign n12175 = n11289 ^ n11288 ;
  assign n12171 = n11433 ^ n11408 ;
  assign n12170 = n12079 ^ n11433 ;
  assign n12172 = n12171 ^ n12170 ;
  assign n12173 = n12084 & ~n12172 ;
  assign n12174 = n12173 ^ n12171 ;
  assign n12176 = n12175 ^ n12174 ;
  assign n12177 = n12176 ^ n11433 ;
  assign n12178 = n10700 & ~n12177 ;
  assign n12179 = n12178 ^ n11433 ;
  assign n12165 = n12086 ^ n12077 ;
  assign n12166 = n12086 ^ n10158 ;
  assign n12167 = n12165 & n12166 ;
  assign n12168 = n12167 ^ n10158 ;
  assign n12169 = n12168 ^ n10179 ;
  assign n12180 = n12179 ^ n12169 ;
  assign n12182 = n12180 ^ x378 ;
  assign n12181 = n12180 ^ n12087 ;
  assign n12183 = n12182 ^ n12181 ;
  assign n12184 = n12092 & ~n12183 ;
  assign n12185 = n12184 ^ n12182 ;
  assign n12186 = n12185 ^ x377 ;
  assign n12188 = n12187 ^ n12186 ;
  assign n12095 = n12072 ^ n12016 ;
  assign n12096 = n12095 ^ n11648 ;
  assign n12097 = n12071 ^ n12070 ;
  assign n12098 = n12097 ^ n11705 ;
  assign n12100 = n11500 ^ n10892 ;
  assign n12101 = n12100 ^ n11522 ;
  assign n12099 = n12069 ^ n12068 ;
  assign n12102 = n12101 ^ n12099 ;
  assign n12104 = n11497 ^ n10885 ;
  assign n12105 = n12104 ^ n11458 ;
  assign n12103 = n12067 ^ n12066 ;
  assign n12106 = n12105 ^ n12103 ;
  assign n12108 = n11494 ^ n11461 ;
  assign n12109 = n12108 ^ n11460 ;
  assign n12107 = n12065 ^ n12063 ;
  assign n12110 = n12109 ^ n12107 ;
  assign n12112 = n11491 ^ n10840 ;
  assign n12113 = n12112 ^ n11463 ;
  assign n12111 = n12062 ^ n12061 ;
  assign n12114 = n12113 ^ n12111 ;
  assign n12116 = n11489 ^ n11466 ;
  assign n12115 = n12060 ^ n12059 ;
  assign n12117 = n12116 ^ n12115 ;
  assign n12119 = n11485 ^ n11470 ;
  assign n12120 = n12119 ^ n11468 ;
  assign n12118 = n12058 ^ n12057 ;
  assign n12121 = n12120 ^ n12118 ;
  assign n12123 = n11483 ^ n11473 ;
  assign n12122 = n12056 ^ n12055 ;
  assign n12124 = n12123 ^ n12122 ;
  assign n12128 = n11479 ^ n11478 ;
  assign n12125 = n11475 ^ n11293 ;
  assign n12126 = n12052 ^ n12051 ;
  assign n12127 = ~n12125 & ~n12126 ;
  assign n12129 = n12128 ^ n12127 ;
  assign n12130 = n12054 ^ n12053 ;
  assign n12131 = n12130 ^ n12127 ;
  assign n12132 = n12129 & ~n12131 ;
  assign n12133 = n12132 ^ n12128 ;
  assign n12134 = n12133 ^ n12122 ;
  assign n12135 = n12124 & n12134 ;
  assign n12136 = n12135 ^ n12123 ;
  assign n12137 = n12136 ^ n12118 ;
  assign n12138 = ~n12121 & ~n12137 ;
  assign n12139 = n12138 ^ n12120 ;
  assign n12140 = n12139 ^ n12115 ;
  assign n12141 = ~n12117 & ~n12140 ;
  assign n12142 = n12141 ^ n12116 ;
  assign n12143 = n12142 ^ n12111 ;
  assign n12144 = ~n12114 & n12143 ;
  assign n12145 = n12144 ^ n12113 ;
  assign n12146 = n12145 ^ n12107 ;
  assign n12147 = n12110 & n12146 ;
  assign n12148 = n12147 ^ n12109 ;
  assign n12149 = n12148 ^ n12103 ;
  assign n12150 = n12106 & ~n12149 ;
  assign n12151 = n12150 ^ n12105 ;
  assign n12152 = n12151 ^ n12099 ;
  assign n12153 = ~n12102 & n12152 ;
  assign n12154 = n12153 ^ n12101 ;
  assign n12155 = n12154 ^ n12097 ;
  assign n12156 = n12098 & n12155 ;
  assign n12157 = n12156 ^ n11705 ;
  assign n12158 = n12157 ^ n12095 ;
  assign n12159 = ~n12096 & ~n12158 ;
  assign n12160 = n12159 ^ n11648 ;
  assign n12094 = n12093 ^ n12073 ;
  assign n12161 = n12160 ^ n12094 ;
  assign n12162 = n12160 ^ n11643 ;
  assign n12163 = ~n12161 & ~n12162 ;
  assign n12164 = n12163 ^ n11643 ;
  assign n12189 = n12188 ^ n12164 ;
  assign n12190 = n12188 ^ n11638 ;
  assign n12191 = n12189 & ~n12190 ;
  assign n12192 = n12191 ^ n11638 ;
  assign n12193 = n12192 ^ n11633 ;
  assign n12212 = n12187 ^ n12180 ;
  assign n12213 = n12185 & ~n12212 ;
  assign n12210 = n12187 ^ n12185 ;
  assign n12211 = ~x377 & n12210 ;
  assign n12214 = n12213 ^ n12211 ;
  assign n12204 = n12175 ^ n11433 ;
  assign n12205 = n12174 & n12204 ;
  assign n12201 = n11291 ^ n11290 ;
  assign n12202 = n12201 ^ n11509 ;
  assign n12203 = n12202 ^ n12175 ;
  assign n12206 = n12205 ^ n12203 ;
  assign n12207 = n12206 ^ n11509 ;
  assign n12208 = n10785 & n12207 ;
  assign n12198 = n11509 ^ n10229 ;
  assign n12197 = n10179 ^ x376 ;
  assign n12199 = n12198 ^ n12197 ;
  assign n12194 = n12179 ^ n12168 ;
  assign n12195 = n12179 ^ n10179 ;
  assign n12196 = n12194 & ~n12195 ;
  assign n12200 = n12199 ^ n12196 ;
  assign n12209 = n12208 ^ n12200 ;
  assign n12215 = n12214 ^ n12209 ;
  assign n12216 = n12215 ^ n12192 ;
  assign n12217 = ~n12193 & ~n12216 ;
  assign n12218 = n12217 ^ n11633 ;
  assign n12233 = n12218 ^ n11297 ;
  assign n12234 = n12231 ^ n11556 ;
  assign n12235 = n12234 ^ n12231 ;
  assign n12236 = n12235 ^ n12218 ;
  assign n12237 = ~n12233 & ~n12236 ;
  assign n12238 = n12237 ^ n12234 ;
  assign n12239 = ~n12232 & ~n12238 ;
  assign n12242 = n12241 ^ n12239 ;
  assign n12244 = n11568 ^ n11559 ;
  assign n12243 = n12240 ^ n12228 ;
  assign n12245 = n12244 ^ n12243 ;
  assign n12246 = n12245 ^ n12228 ;
  assign n12247 = n12242 & ~n12246 ;
  assign n12248 = n12247 ^ n12243 ;
  assign n12249 = ~n12229 & ~n12248 ;
  assign n12251 = n12250 ^ n12249 ;
  assign n12252 = ~n12226 & n12251 ;
  assign n12224 = n11624 ^ n11619 ;
  assign n12253 = n12252 ^ n12224 ;
  assign n12254 = n12025 ^ n12024 ;
  assign n12255 = n12254 ^ n11619 ;
  assign n12256 = ~n12253 & n12255 ;
  assign n12223 = n11619 ^ n11614 ;
  assign n12257 = n12256 ^ n12223 ;
  assign n12258 = n12027 ^ n12026 ;
  assign n12259 = n12258 ^ n11614 ;
  assign n12260 = ~n12257 & ~n12259 ;
  assign n12222 = n11614 ^ n11609 ;
  assign n12261 = n12260 ^ n12222 ;
  assign n12262 = n12029 ^ n12028 ;
  assign n12263 = n12262 ^ n11609 ;
  assign n12264 = n12261 & n12263 ;
  assign n12221 = n11609 ^ n11604 ;
  assign n12265 = n12264 ^ n12221 ;
  assign n12220 = n12031 ^ n12030 ;
  assign n12416 = n12220 ^ n11604 ;
  assign n12417 = n12265 & n12416 ;
  assign n12419 = n12418 ^ n12417 ;
  assign n12415 = n12033 ^ n12032 ;
  assign n12580 = n12415 ^ n11768 ;
  assign n12581 = n12419 & n12580 ;
  assign n12582 = n12581 ^ n11768 ;
  assign n12579 = n12035 ^ n12034 ;
  assign n12583 = n12582 ^ n12579 ;
  assign n12597 = n12582 ^ n11779 ;
  assign n12598 = ~n12583 & n12597 ;
  assign n12599 = n12598 ^ n11779 ;
  assign n12665 = n12664 ^ n12599 ;
  assign n12600 = n12037 ^ n12036 ;
  assign n12666 = n12664 ^ n12600 ;
  assign n12667 = ~n12665 & n12666 ;
  assign n12663 = n12600 ^ n11966 ;
  assign n12668 = n12667 ^ n12663 ;
  assign n12784 = n11986 ^ n11370 ;
  assign n12785 = n12784 ^ n11966 ;
  assign n12669 = n12039 ^ n12038 ;
  assign n12786 = n12785 ^ n12669 ;
  assign n12787 = n12786 ^ n12784 ;
  assign n12788 = ~n12668 & n12787 ;
  assign n12789 = n12788 ^ n12785 ;
  assign n12790 = n12041 ^ n12040 ;
  assign n12817 = n12790 ^ n12784 ;
  assign n12818 = n12789 & ~n12817 ;
  assign n12816 = n12784 ^ n12006 ;
  assign n12819 = n12818 ^ n12816 ;
  assign n12833 = n12084 ^ n11408 ;
  assign n12834 = n12833 ^ n12006 ;
  assign n12815 = n12043 ^ n12042 ;
  assign n12835 = n12834 ^ n12815 ;
  assign n12836 = n12835 ^ n12833 ;
  assign n12837 = ~n12819 & ~n12836 ;
  assign n12838 = n12837 ^ n12834 ;
  assign n12839 = n12045 ^ n12044 ;
  assign n12864 = n12839 ^ n12833 ;
  assign n12865 = n12838 & ~n12864 ;
  assign n12863 = n12833 ^ n12176 ;
  assign n12866 = n12865 ^ n12863 ;
  assign n12862 = n12048 ^ n12046 ;
  assign n12915 = n12862 ^ n12176 ;
  assign n12916 = n12866 & n12915 ;
  assign n12913 = n12050 ^ n12049 ;
  assign n12912 = n12862 ^ n12206 ;
  assign n12914 = n12913 ^ n12912 ;
  assign n12917 = n12916 ^ n12914 ;
  assign n12918 = n12917 ^ n12206 ;
  assign n12919 = ~n11509 & n12918 ;
  assign n12909 = n12206 ^ n10785 ;
  assign n12908 = n10700 ^ x24 ;
  assign n12910 = n12909 ^ n12908 ;
  assign n12867 = n12866 ^ n12862 ;
  assign n12868 = n12867 ^ n12176 ;
  assign n12869 = ~n11433 & ~n12868 ;
  assign n12870 = n12869 ^ n12176 ;
  assign n12820 = n12819 ^ n12815 ;
  assign n12821 = n12820 ^ n12006 ;
  assign n12822 = n11391 & n12821 ;
  assign n12823 = n12822 ^ n12006 ;
  assign n12601 = n12600 ^ n12599 ;
  assign n12602 = n11331 & ~n12601 ;
  assign n12603 = n12602 ^ n11949 ;
  assign n12420 = n12419 ^ n12415 ;
  assign n12421 = n12420 ^ n11768 ;
  assign n12422 = n11242 & n12421 ;
  assign n12423 = n12422 ^ n11768 ;
  assign n12266 = n12265 ^ n12220 ;
  assign n12267 = n12266 ^ n11604 ;
  assign n12268 = ~n11227 & n12267 ;
  assign n12269 = n12268 ^ n11604 ;
  assign n12270 = n12269 ^ n11220 ;
  assign n12271 = n12262 ^ n12261 ;
  assign n12272 = n12271 ^ n11609 ;
  assign n12273 = n11204 & n12272 ;
  assign n12274 = n12273 ^ n11609 ;
  assign n12275 = n12274 ^ n11197 ;
  assign n12276 = n12258 ^ n12257 ;
  assign n12277 = n12276 ^ n11614 ;
  assign n12278 = ~n11181 & n12277 ;
  assign n12279 = n12278 ^ n11614 ;
  assign n12280 = n12279 ^ n11174 ;
  assign n12281 = n12254 ^ n12253 ;
  assign n12282 = n12281 ^ n11619 ;
  assign n12283 = n11158 & ~n12282 ;
  assign n12284 = n12283 ^ n11619 ;
  assign n12285 = n12284 ^ n11151 ;
  assign n12286 = n12251 ^ n12225 ;
  assign n12287 = n12286 ^ n11624 ;
  assign n12288 = n11133 & ~n12287 ;
  assign n12289 = n12288 ^ n11624 ;
  assign n12290 = n12289 ^ n11130 ;
  assign n12291 = ~n11573 & n12248 ;
  assign n12292 = n12291 ^ n11572 ;
  assign n12293 = n12292 ^ n11127 ;
  assign n12294 = n11559 & ~n12242 ;
  assign n12295 = n12294 ^ n11568 ;
  assign n12296 = n12295 ^ n11003 ;
  assign n12384 = n12238 ^ n12230 ;
  assign n12385 = n12384 ^ n12231 ;
  assign n12386 = ~n10988 & n12385 ;
  assign n12387 = n12386 ^ n12231 ;
  assign n12301 = ~n10941 & ~n12189 ;
  assign n12302 = n12301 ^ n11638 ;
  assign n12303 = n12302 ^ n10934 ;
  assign n12367 = ~n10925 & n12161 ;
  assign n12368 = n12367 ^ n11643 ;
  assign n12361 = n10910 & n12158 ;
  assign n12362 = n12361 ^ n11648 ;
  assign n12304 = n11298 & ~n12155 ;
  assign n12305 = n12304 ^ n11705 ;
  assign n12306 = n12305 ^ n10837 ;
  assign n12307 = ~n10892 & ~n12152 ;
  assign n12308 = n12307 ^ n12101 ;
  assign n12309 = n12308 ^ n9886 ;
  assign n12349 = n10885 & n12149 ;
  assign n12350 = n12349 ^ n12105 ;
  assign n12310 = n11461 & ~n12146 ;
  assign n12311 = n12310 ^ n12109 ;
  assign n12312 = n12311 ^ n10822 ;
  assign n12313 = ~n10840 & ~n12143 ;
  assign n12314 = n12313 ^ n12113 ;
  assign n12315 = n12314 ^ n9934 ;
  assign n12316 = n11465 & n12140 ;
  assign n12317 = n12316 ^ n12116 ;
  assign n12318 = n12317 ^ n9938 ;
  assign n12319 = n11470 & n12137 ;
  assign n12320 = n12319 ^ n12120 ;
  assign n12321 = n12320 ^ n10794 ;
  assign n12322 = n11472 & ~n12134 ;
  assign n12323 = n12322 ^ n12123 ;
  assign n12324 = n12323 ^ n10797 ;
  assign n12325 = n11475 & n12126 ;
  assign n12326 = n12325 ^ n11293 ;
  assign n12327 = n9533 & ~n12326 ;
  assign n12328 = n12327 ^ n10803 ;
  assign n12329 = n11477 & n12131 ;
  assign n12330 = n12329 ^ n12128 ;
  assign n12331 = n12330 ^ n12327 ;
  assign n12332 = n12328 & ~n12331 ;
  assign n12333 = n12332 ^ n10803 ;
  assign n12334 = n12333 ^ n12323 ;
  assign n12335 = ~n12324 & n12334 ;
  assign n12336 = n12335 ^ n10797 ;
  assign n12337 = n12336 ^ n12320 ;
  assign n12338 = n12321 & ~n12337 ;
  assign n12339 = n12338 ^ n10794 ;
  assign n12340 = n12339 ^ n12317 ;
  assign n12341 = n12318 & n12340 ;
  assign n12342 = n12341 ^ n9938 ;
  assign n12343 = n12342 ^ n12314 ;
  assign n12344 = ~n12315 & ~n12343 ;
  assign n12345 = n12344 ^ n9934 ;
  assign n12346 = n12345 ^ n12311 ;
  assign n12347 = n12312 & ~n12346 ;
  assign n12348 = n12347 ^ n10822 ;
  assign n12351 = n12350 ^ n12348 ;
  assign n12352 = n12350 ^ n9930 ;
  assign n12353 = ~n12351 & n12352 ;
  assign n12354 = n12353 ^ n9930 ;
  assign n12355 = n12354 ^ n12308 ;
  assign n12356 = ~n12309 & ~n12355 ;
  assign n12357 = n12356 ^ n9886 ;
  assign n12358 = n12357 ^ n12305 ;
  assign n12359 = ~n12306 & ~n12358 ;
  assign n12360 = n12359 ^ n10837 ;
  assign n12363 = n12362 ^ n12360 ;
  assign n12364 = n12362 ^ n10907 ;
  assign n12365 = ~n12363 & n12364 ;
  assign n12366 = n12365 ^ n10907 ;
  assign n12369 = n12368 ^ n12366 ;
  assign n12370 = n12368 ^ n10918 ;
  assign n12371 = n12369 & ~n12370 ;
  assign n12372 = n12371 ^ n10918 ;
  assign n12373 = n12372 ^ n12302 ;
  assign n12374 = n12303 & n12373 ;
  assign n12375 = n12374 ^ n10934 ;
  assign n12299 = n10957 & n12216 ;
  assign n12300 = n12299 ^ n11633 ;
  assign n12376 = n12375 ^ n12300 ;
  assign n12377 = n12375 ^ n10950 ;
  assign n12378 = n12376 & ~n12377 ;
  assign n12379 = n12378 ^ n10950 ;
  assign n12297 = ~n10973 & n12233 ;
  assign n12298 = n12297 ^ n11556 ;
  assign n12380 = n12379 ^ n12298 ;
  assign n12381 = n12379 ^ n10966 ;
  assign n12382 = n12380 & n12381 ;
  assign n12383 = n12382 ^ n10966 ;
  assign n12388 = n12387 ^ n12383 ;
  assign n12389 = n12295 ^ n10981 ;
  assign n12390 = n12389 ^ n12295 ;
  assign n12391 = n12390 ^ n12383 ;
  assign n12392 = ~n12388 & ~n12391 ;
  assign n12393 = n12392 ^ n12389 ;
  assign n12394 = n12296 & ~n12393 ;
  assign n12395 = n12394 ^ n11003 ;
  assign n12396 = n12395 ^ n12292 ;
  assign n12397 = n12293 & ~n12396 ;
  assign n12398 = n12397 ^ n11127 ;
  assign n12399 = n12398 ^ n12289 ;
  assign n12400 = ~n12290 & ~n12399 ;
  assign n12401 = n12400 ^ n11130 ;
  assign n12402 = n12401 ^ n12284 ;
  assign n12403 = ~n12285 & ~n12402 ;
  assign n12404 = n12403 ^ n11151 ;
  assign n12405 = n12404 ^ n12279 ;
  assign n12406 = ~n12280 & ~n12405 ;
  assign n12407 = n12406 ^ n11174 ;
  assign n12408 = n12407 ^ n12274 ;
  assign n12409 = ~n12275 & n12408 ;
  assign n12410 = n12409 ^ n11197 ;
  assign n12411 = n12410 ^ n12269 ;
  assign n12412 = n12270 & n12411 ;
  assign n12413 = n12412 ^ n11220 ;
  assign n12578 = n12423 ^ n12413 ;
  assign n12584 = ~n11775 & n12583 ;
  assign n12585 = n12584 ^ n11779 ;
  assign n12586 = n12585 ^ n10450 ;
  assign n12587 = n12586 ^ n12413 ;
  assign n12588 = n12587 ^ n12585 ;
  assign n12589 = ~n12578 & ~n12588 ;
  assign n12590 = n12589 ^ n12586 ;
  assign n12593 = n12585 ^ n10324 ;
  assign n12594 = n12590 & n12593 ;
  assign n12595 = n12594 ^ n10324 ;
  assign n12662 = n12603 ^ n12595 ;
  assign n12670 = n12669 ^ n12668 ;
  assign n12671 = n12670 ^ n11966 ;
  assign n12672 = n11959 & ~n12671 ;
  assign n12673 = n12672 ^ n11966 ;
  assign n12674 = n12673 ^ n11324 ;
  assign n12675 = n12674 ^ n12595 ;
  assign n12676 = n12675 ^ n12673 ;
  assign n12677 = ~n12662 & ~n12676 ;
  assign n12678 = n12677 ^ n12674 ;
  assign n12795 = n12673 ^ n10622 ;
  assign n12796 = ~n12678 & ~n12795 ;
  assign n12797 = n12796 ^ n10622 ;
  assign n12798 = n12797 ^ n10635 ;
  assign n12791 = n12790 ^ n12789 ;
  assign n12792 = n12791 ^ n11986 ;
  assign n12793 = ~n11370 & ~n12792 ;
  assign n12794 = n12793 ^ n12791 ;
  assign n12811 = n12797 ^ n12794 ;
  assign n12812 = ~n12798 & ~n12811 ;
  assign n12813 = n12812 ^ n10635 ;
  assign n12844 = n12823 ^ n12813 ;
  assign n12845 = n12823 ^ n10660 ;
  assign n12846 = n12844 & ~n12845 ;
  assign n12847 = n12846 ^ n10660 ;
  assign n12840 = n12839 ^ n12838 ;
  assign n12841 = n12840 ^ n12084 ;
  assign n12842 = ~n11408 & ~n12841 ;
  assign n12843 = n12842 ^ n12840 ;
  assign n12857 = n12847 ^ n12843 ;
  assign n12858 = n12843 ^ n11401 ;
  assign n12859 = ~n12857 & ~n12858 ;
  assign n12860 = n12859 ^ n11401 ;
  assign n12905 = n12870 ^ n12860 ;
  assign n12906 = n12870 ^ n10700 ;
  assign n12907 = n12905 & n12906 ;
  assign n12911 = n12910 ^ n12907 ;
  assign n12920 = n12919 ^ n12911 ;
  assign n12591 = n12590 ^ n10324 ;
  assign n12414 = n12413 ^ n10450 ;
  assign n12424 = n12423 ^ n12414 ;
  assign n12425 = n12424 ^ x16 ;
  assign n12427 = n12381 ^ n12298 ;
  assign n12428 = n12427 ^ x9 ;
  assign n12506 = n12372 ^ n10934 ;
  assign n12507 = n12506 ^ n12302 ;
  assign n12429 = n12366 ^ n10918 ;
  assign n12430 = n12429 ^ n12368 ;
  assign n12431 = n12430 ^ x12 ;
  assign n12433 = n12326 ^ n9533 ;
  assign n12434 = x7 & ~n12433 ;
  assign n12432 = n12330 ^ n12328 ;
  assign n12435 = n12434 ^ n12432 ;
  assign n12436 = n12333 ^ n10797 ;
  assign n12437 = n12436 ^ n12323 ;
  assign n12438 = n12437 ^ x6 ;
  assign n12439 = n12438 ^ n12432 ;
  assign n12440 = n12439 ^ n12437 ;
  assign n12441 = ~n12435 & n12440 ;
  assign n12442 = n12441 ^ n12438 ;
  assign n12443 = n12336 ^ n10794 ;
  assign n12444 = n12443 ^ n12320 ;
  assign n12446 = n12444 ^ x5 ;
  assign n12445 = n12444 ^ n12437 ;
  assign n12447 = n12446 ^ n12445 ;
  assign n12448 = n12442 & ~n12447 ;
  assign n12449 = n12448 ^ n12446 ;
  assign n12450 = n12339 ^ n9938 ;
  assign n12451 = n12450 ^ n12317 ;
  assign n12453 = n12451 ^ x4 ;
  assign n12452 = n12451 ^ n12444 ;
  assign n12454 = n12453 ^ n12452 ;
  assign n12455 = ~n12449 & n12454 ;
  assign n12456 = n12455 ^ n12453 ;
  assign n12457 = n12342 ^ n9934 ;
  assign n12458 = n12457 ^ n12314 ;
  assign n12460 = n12458 ^ x3 ;
  assign n12459 = n12458 ^ n12451 ;
  assign n12461 = n12460 ^ n12459 ;
  assign n12462 = ~n12456 & n12461 ;
  assign n12463 = n12462 ^ n12460 ;
  assign n12464 = n12345 ^ n10822 ;
  assign n12465 = n12464 ^ n12311 ;
  assign n12467 = n12465 ^ x2 ;
  assign n12466 = n12465 ^ n12458 ;
  assign n12468 = n12467 ^ n12466 ;
  assign n12469 = ~n12463 & n12468 ;
  assign n12470 = n12469 ^ n12467 ;
  assign n12471 = n12348 ^ n9930 ;
  assign n12472 = n12471 ^ n12350 ;
  assign n12474 = n12472 ^ x1 ;
  assign n12473 = n12472 ^ n12465 ;
  assign n12475 = n12474 ^ n12473 ;
  assign n12476 = ~n12470 & n12475 ;
  assign n12477 = n12476 ^ n12474 ;
  assign n12478 = n12354 ^ n9886 ;
  assign n12479 = n12478 ^ n12308 ;
  assign n12481 = n12479 ^ x0 ;
  assign n12480 = n12479 ^ n12472 ;
  assign n12482 = n12481 ^ n12480 ;
  assign n12483 = ~n12477 & n12482 ;
  assign n12484 = n12483 ^ n12481 ;
  assign n12485 = n12357 ^ n10837 ;
  assign n12486 = n12485 ^ n12305 ;
  assign n12488 = n12486 ^ x15 ;
  assign n12487 = n12486 ^ n12479 ;
  assign n12489 = n12488 ^ n12487 ;
  assign n12490 = n12484 & ~n12489 ;
  assign n12491 = n12490 ^ n12488 ;
  assign n12492 = n12360 ^ n10907 ;
  assign n12493 = n12492 ^ n12362 ;
  assign n12495 = n12493 ^ x14 ;
  assign n12494 = n12493 ^ n12486 ;
  assign n12496 = n12495 ^ n12494 ;
  assign n12497 = ~n12491 & n12496 ;
  assign n12498 = n12497 ^ n12495 ;
  assign n12500 = n12430 ^ x13 ;
  assign n12499 = n12493 ^ n12430 ;
  assign n12501 = n12500 ^ n12499 ;
  assign n12502 = ~n12498 & n12501 ;
  assign n12503 = n12502 ^ n12500 ;
  assign n12504 = ~n12431 & n12503 ;
  assign n12505 = n12504 ^ x12 ;
  assign n12508 = n12507 ^ n12505 ;
  assign n12509 = n12377 ^ n12300 ;
  assign n12510 = n12509 ^ x11 ;
  assign n12511 = n12510 ^ n12505 ;
  assign n12512 = n12511 ^ n12509 ;
  assign n12513 = ~n12508 & n12512 ;
  assign n12514 = n12513 ^ n12510 ;
  assign n12516 = n12427 ^ x10 ;
  assign n12515 = n12509 ^ n12427 ;
  assign n12517 = n12516 ^ n12515 ;
  assign n12518 = n12514 & ~n12517 ;
  assign n12519 = n12518 ^ n12516 ;
  assign n12520 = ~n12428 & n12519 ;
  assign n12521 = n12520 ^ x9 ;
  assign n12522 = n12521 ^ x8 ;
  assign n12523 = n12383 ^ n10981 ;
  assign n12524 = n12523 ^ n12387 ;
  assign n12525 = n12524 ^ n12521 ;
  assign n12526 = n12522 & n12525 ;
  assign n12527 = n12526 ^ x8 ;
  assign n12426 = n12393 ^ n11003 ;
  assign n12528 = n12527 ^ n12426 ;
  assign n12529 = n12395 ^ n11127 ;
  assign n12530 = n12529 ^ n12292 ;
  assign n12531 = n12530 ^ x23 ;
  assign n12532 = n12531 ^ n12426 ;
  assign n12533 = n12532 ^ n12530 ;
  assign n12534 = n12528 & ~n12533 ;
  assign n12535 = n12534 ^ n12531 ;
  assign n12536 = n12398 ^ n11130 ;
  assign n12537 = n12536 ^ n12289 ;
  assign n12539 = n12537 ^ x22 ;
  assign n12538 = n12537 ^ n12530 ;
  assign n12540 = n12539 ^ n12538 ;
  assign n12541 = n12535 & ~n12540 ;
  assign n12542 = n12541 ^ n12539 ;
  assign n12543 = n12401 ^ n11151 ;
  assign n12544 = n12543 ^ n12284 ;
  assign n12546 = n12544 ^ x21 ;
  assign n12545 = n12544 ^ n12537 ;
  assign n12547 = n12546 ^ n12545 ;
  assign n12548 = ~n12542 & n12547 ;
  assign n12549 = n12548 ^ n12546 ;
  assign n12550 = n12404 ^ n11174 ;
  assign n12551 = n12550 ^ n12279 ;
  assign n12553 = n12551 ^ x20 ;
  assign n12552 = n12551 ^ n12544 ;
  assign n12554 = n12553 ^ n12552 ;
  assign n12555 = n12549 & ~n12554 ;
  assign n12556 = n12555 ^ n12553 ;
  assign n12557 = n12407 ^ n11197 ;
  assign n12558 = n12557 ^ n12274 ;
  assign n12560 = n12558 ^ x19 ;
  assign n12559 = n12558 ^ n12551 ;
  assign n12561 = n12560 ^ n12559 ;
  assign n12562 = ~n12556 & n12561 ;
  assign n12563 = n12562 ^ n12560 ;
  assign n12564 = n12410 ^ n11220 ;
  assign n12565 = n12564 ^ n12269 ;
  assign n12567 = n12565 ^ x18 ;
  assign n12566 = n12565 ^ n12558 ;
  assign n12568 = n12567 ^ n12566 ;
  assign n12569 = n12563 & ~n12568 ;
  assign n12570 = n12569 ^ n12567 ;
  assign n12572 = n12424 ^ x17 ;
  assign n12571 = n12565 ^ n12424 ;
  assign n12573 = n12572 ^ n12571 ;
  assign n12574 = ~n12570 & n12573 ;
  assign n12575 = n12574 ^ n12572 ;
  assign n12576 = n12425 & ~n12575 ;
  assign n12577 = n12576 ^ x16 ;
  assign n12592 = n12591 ^ n12577 ;
  assign n12596 = n12595 ^ n11324 ;
  assign n12604 = n12603 ^ n12596 ;
  assign n12605 = n12604 ^ x31 ;
  assign n12606 = n12605 ^ n12577 ;
  assign n12607 = n12606 ^ n12604 ;
  assign n12608 = ~n12592 & n12607 ;
  assign n12609 = n12608 ^ n12605 ;
  assign n12679 = n12678 ^ n10622 ;
  assign n12681 = n12679 ^ x30 ;
  assign n12680 = n12679 ^ n12604 ;
  assign n12682 = n12681 ^ n12680 ;
  assign n12683 = ~n12609 & n12682 ;
  assign n12684 = n12683 ^ n12681 ;
  assign n12799 = n12798 ^ n12794 ;
  assign n12801 = n12799 ^ x29 ;
  assign n12800 = n12799 ^ n12679 ;
  assign n12802 = n12801 ^ n12800 ;
  assign n12803 = n12684 & ~n12802 ;
  assign n12804 = n12803 ^ n12801 ;
  assign n12814 = n12813 ^ n10660 ;
  assign n12824 = n12823 ^ n12814 ;
  assign n12826 = n12824 ^ x28 ;
  assign n12825 = n12824 ^ n12799 ;
  assign n12827 = n12826 ^ n12825 ;
  assign n12828 = ~n12804 & n12827 ;
  assign n12829 = n12828 ^ n12826 ;
  assign n12848 = n12847 ^ n11401 ;
  assign n12849 = n12848 ^ n12843 ;
  assign n12851 = n12849 ^ x27 ;
  assign n12850 = n12849 ^ n12824 ;
  assign n12852 = n12851 ^ n12850 ;
  assign n12853 = n12829 & ~n12852 ;
  assign n12854 = n12853 ^ n12851 ;
  assign n12861 = n12860 ^ n10700 ;
  assign n12871 = n12870 ^ n12861 ;
  assign n12873 = n12871 ^ x26 ;
  assign n12872 = n12871 ^ n12849 ;
  assign n12874 = n12873 ^ n12872 ;
  assign n12875 = n12854 & ~n12874 ;
  assign n12876 = n12875 ^ n12873 ;
  assign n12830 = n12829 ^ x27 ;
  assign n12610 = n12609 ^ x30 ;
  assign n12611 = n12508 ^ x11 ;
  assign n12612 = n12434 ^ x6 ;
  assign n12613 = n12612 ^ n12432 ;
  assign n12614 = n12442 ^ x5 ;
  assign n12615 = n12613 & ~n12614 ;
  assign n12616 = n12449 ^ x4 ;
  assign n12617 = ~n12615 & ~n12616 ;
  assign n12618 = n12456 ^ x3 ;
  assign n12619 = ~n12617 & n12618 ;
  assign n12620 = n12463 ^ x2 ;
  assign n12621 = ~n12619 & ~n12620 ;
  assign n12622 = n12470 ^ x1 ;
  assign n12623 = ~n12621 & n12622 ;
  assign n12624 = n12477 ^ x0 ;
  assign n12625 = ~n12623 & ~n12624 ;
  assign n12626 = n12484 ^ x15 ;
  assign n12627 = n12625 & n12626 ;
  assign n12628 = n12491 ^ x14 ;
  assign n12629 = n12627 & ~n12628 ;
  assign n12630 = n12498 ^ x13 ;
  assign n12631 = n12629 & ~n12630 ;
  assign n12632 = n12503 ^ x12 ;
  assign n12633 = ~n12631 & ~n12632 ;
  assign n12634 = n12611 & n12633 ;
  assign n12635 = n12514 ^ x10 ;
  assign n12636 = n12634 & ~n12635 ;
  assign n12637 = n12519 ^ x9 ;
  assign n12638 = ~n12636 & n12637 ;
  assign n12639 = n12525 ^ x8 ;
  assign n12640 = n12638 & n12639 ;
  assign n12641 = n12527 ^ x23 ;
  assign n12642 = n12641 ^ n12426 ;
  assign n12643 = ~n12640 & ~n12642 ;
  assign n12644 = n12535 ^ x22 ;
  assign n12645 = ~n12643 & n12644 ;
  assign n12646 = n12542 ^ x21 ;
  assign n12647 = n12645 & ~n12646 ;
  assign n12648 = n12549 ^ x20 ;
  assign n12649 = ~n12647 & ~n12648 ;
  assign n12650 = n12556 ^ x19 ;
  assign n12651 = ~n12649 & ~n12650 ;
  assign n12652 = n12563 ^ x18 ;
  assign n12653 = n12651 & n12652 ;
  assign n12654 = n12570 ^ x17 ;
  assign n12655 = ~n12653 & n12654 ;
  assign n12656 = n12575 ^ x16 ;
  assign n12657 = ~n12655 & ~n12656 ;
  assign n12658 = n12577 ^ x31 ;
  assign n12659 = n12658 ^ n12591 ;
  assign n12660 = n12657 & ~n12659 ;
  assign n12661 = n12610 & ~n12660 ;
  assign n12685 = n12684 ^ x29 ;
  assign n12783 = n12661 & ~n12685 ;
  assign n12805 = n12804 ^ x28 ;
  assign n12831 = ~n12783 & ~n12805 ;
  assign n12832 = ~n12830 & ~n12831 ;
  assign n12855 = n12854 ^ x26 ;
  assign n12856 = ~n12832 & n12855 ;
  assign n12900 = n12871 ^ n12856 ;
  assign n12903 = n12876 & ~n12900 ;
  assign n12899 = n12876 ^ n12871 ;
  assign n12901 = n12900 ^ n12899 ;
  assign n12902 = x25 & ~n12901 ;
  assign n12904 = n12903 ^ n12902 ;
  assign n12921 = n12920 ^ n12904 ;
  assign n12877 = n12876 ^ x25 ;
  assign n12878 = n12877 ^ n12856 ;
  assign n12879 = n12878 ^ n12286 ;
  assign n12881 = n12248 ^ n12227 ;
  assign n12880 = n12855 ^ n12832 ;
  assign n12882 = n12881 ^ n12880 ;
  assign n12884 = n12244 ^ n12242 ;
  assign n12883 = n12831 ^ n12830 ;
  assign n12885 = n12884 ^ n12883 ;
  assign n12806 = n12805 ^ n12783 ;
  assign n12886 = n12806 ^ n12384 ;
  assign n12686 = n12685 ^ n12661 ;
  assign n11557 = n11556 ^ n11297 ;
  assign n12219 = n12218 ^ n11557 ;
  assign n12687 = n12686 ^ n12219 ;
  assign n12689 = n12215 ^ n12193 ;
  assign n12688 = n12660 ^ n12610 ;
  assign n12690 = n12689 ^ n12688 ;
  assign n12692 = n12164 ^ n11638 ;
  assign n12693 = n12692 ^ n12188 ;
  assign n12691 = n12659 ^ n12657 ;
  assign n12694 = n12693 ^ n12691 ;
  assign n12696 = n12162 ^ n12094 ;
  assign n12772 = n12696 ^ n12691 ;
  assign n12695 = n12656 ^ n12655 ;
  assign n12697 = n12696 ^ n12695 ;
  assign n12699 = n12157 ^ n11648 ;
  assign n12700 = n12699 ^ n12095 ;
  assign n12698 = n12654 ^ n12653 ;
  assign n12701 = n12700 ^ n12698 ;
  assign n12703 = n12154 ^ n11705 ;
  assign n12704 = n12703 ^ n12097 ;
  assign n12702 = n12652 ^ n12651 ;
  assign n12705 = n12704 ^ n12702 ;
  assign n12707 = n12151 ^ n12101 ;
  assign n12708 = n12707 ^ n12099 ;
  assign n12706 = n12650 ^ n12649 ;
  assign n12709 = n12708 ^ n12706 ;
  assign n12711 = n12148 ^ n12105 ;
  assign n12712 = n12711 ^ n12103 ;
  assign n12710 = n12648 ^ n12647 ;
  assign n12713 = n12712 ^ n12710 ;
  assign n12715 = n12145 ^ n12109 ;
  assign n12716 = n12715 ^ n12107 ;
  assign n12714 = n12646 ^ n12645 ;
  assign n12717 = n12716 ^ n12714 ;
  assign n12720 = n12644 ^ n12643 ;
  assign n12718 = n12142 ^ n12113 ;
  assign n12719 = n12718 ^ n12111 ;
  assign n12721 = n12720 ^ n12719 ;
  assign n12723 = n12139 ^ n12116 ;
  assign n12724 = n12723 ^ n12115 ;
  assign n12722 = n12642 ^ n12640 ;
  assign n12725 = n12724 ^ n12722 ;
  assign n12728 = n12639 ^ n12638 ;
  assign n12726 = n12136 ^ n12120 ;
  assign n12727 = n12726 ^ n12118 ;
  assign n12729 = n12728 ^ n12727 ;
  assign n12731 = n12133 ^ n12123 ;
  assign n12732 = n12731 ^ n12122 ;
  assign n12730 = n12637 ^ n12636 ;
  assign n12733 = n12732 ^ n12730 ;
  assign n12737 = n12130 ^ n12129 ;
  assign n12734 = n12633 ^ n12611 ;
  assign n12735 = n12126 ^ n12125 ;
  assign n12736 = n12734 & n12735 ;
  assign n12738 = n12737 ^ n12736 ;
  assign n12739 = n12635 ^ n12634 ;
  assign n12740 = n12739 ^ n12736 ;
  assign n12741 = n12738 & n12740 ;
  assign n12742 = n12741 ^ n12737 ;
  assign n12743 = n12742 ^ n12730 ;
  assign n12744 = n12733 & ~n12743 ;
  assign n12745 = n12744 ^ n12732 ;
  assign n12746 = n12745 ^ n12727 ;
  assign n12747 = ~n12729 & ~n12746 ;
  assign n12748 = n12747 ^ n12728 ;
  assign n12749 = n12748 ^ n12722 ;
  assign n12750 = ~n12725 & n12749 ;
  assign n12751 = n12750 ^ n12724 ;
  assign n12752 = n12751 ^ n12719 ;
  assign n12753 = n12721 & n12752 ;
  assign n12754 = n12753 ^ n12720 ;
  assign n12755 = n12754 ^ n12714 ;
  assign n12756 = ~n12717 & ~n12755 ;
  assign n12757 = n12756 ^ n12716 ;
  assign n12758 = n12757 ^ n12710 ;
  assign n12759 = n12713 & n12758 ;
  assign n12760 = n12759 ^ n12712 ;
  assign n12761 = n12760 ^ n12706 ;
  assign n12762 = n12709 & n12761 ;
  assign n12763 = n12762 ^ n12708 ;
  assign n12764 = n12763 ^ n12702 ;
  assign n12765 = ~n12705 & ~n12764 ;
  assign n12766 = n12765 ^ n12704 ;
  assign n12767 = n12766 ^ n12698 ;
  assign n12768 = ~n12701 & n12767 ;
  assign n12769 = n12768 ^ n12700 ;
  assign n12770 = n12769 ^ n12695 ;
  assign n12771 = n12697 & n12770 ;
  assign n12773 = n12772 ^ n12771 ;
  assign n12774 = n12694 & n12773 ;
  assign n12775 = n12774 ^ n12693 ;
  assign n12776 = n12775 ^ n12688 ;
  assign n12777 = ~n12690 & n12776 ;
  assign n12778 = n12777 ^ n12689 ;
  assign n12779 = n12778 ^ n12219 ;
  assign n12780 = n12687 & n12779 ;
  assign n12781 = n12780 ^ n12686 ;
  assign n12887 = n12806 ^ n12781 ;
  assign n12888 = ~n12886 & ~n12887 ;
  assign n12889 = n12888 ^ n12384 ;
  assign n12890 = n12889 ^ n12883 ;
  assign n12891 = ~n12885 & ~n12890 ;
  assign n12892 = n12891 ^ n12884 ;
  assign n12893 = n12892 ^ n12880 ;
  assign n12894 = ~n12882 & n12893 ;
  assign n12895 = n12894 ^ n12881 ;
  assign n12896 = n12895 ^ n12878 ;
  assign n12897 = ~n12879 & ~n12896 ;
  assign n12898 = n12897 ^ n12286 ;
  assign n12922 = n12921 ^ n12898 ;
  assign n12959 = n11619 & ~n12922 ;
  assign n12960 = n12959 ^ n12281 ;
  assign n12961 = n12960 ^ n11158 ;
  assign n12962 = ~n11624 & n12896 ;
  assign n12963 = n12962 ^ n12286 ;
  assign n12964 = n12963 ^ n11133 ;
  assign n12965 = ~n12244 & ~n12890 ;
  assign n12966 = n12965 ^ n12242 ;
  assign n12967 = n12966 ^ n11559 ;
  assign n13058 = n12231 & n12887 ;
  assign n13059 = n13058 ^ n12384 ;
  assign n12968 = n12778 ^ n12686 ;
  assign n12969 = ~n11556 & ~n12968 ;
  assign n12970 = n12969 ^ n12219 ;
  assign n12971 = n12970 ^ n10973 ;
  assign n12972 = n11633 & ~n12776 ;
  assign n12973 = n12972 ^ n12689 ;
  assign n12974 = n12973 ^ n10957 ;
  assign n12975 = n11648 & ~n12767 ;
  assign n12976 = n12975 ^ n12700 ;
  assign n12977 = n12976 ^ n10910 ;
  assign n12978 = ~n11705 & n12764 ;
  assign n12979 = n12978 ^ n12704 ;
  assign n12980 = n12979 ^ n11298 ;
  assign n12981 = n12101 & ~n12761 ;
  assign n12982 = n12981 ^ n12708 ;
  assign n12983 = n12982 ^ n10892 ;
  assign n12984 = n12105 & ~n12758 ;
  assign n12985 = n12984 ^ n12712 ;
  assign n12986 = n12985 ^ n10885 ;
  assign n12987 = ~n12123 & n12743 ;
  assign n12988 = n12987 ^ n12732 ;
  assign n12989 = n12988 ^ n11472 ;
  assign n12990 = ~n12125 & ~n12734 ;
  assign n12991 = n12990 ^ n12126 ;
  assign n12992 = n11475 & ~n12991 ;
  assign n12993 = n12992 ^ n11477 ;
  assign n12995 = n12128 & ~n12740 ;
  assign n12994 = n12992 ^ n12737 ;
  assign n12996 = n12995 ^ n12994 ;
  assign n12997 = n12993 & ~n12996 ;
  assign n12998 = n12997 ^ n11477 ;
  assign n12999 = n12998 ^ n12988 ;
  assign n13000 = n12989 & ~n12999 ;
  assign n13001 = n13000 ^ n11472 ;
  assign n13002 = n13001 ^ n11470 ;
  assign n13003 = n12745 ^ n12728 ;
  assign n13004 = n12120 & ~n13003 ;
  assign n13005 = n13004 ^ n12727 ;
  assign n13006 = n13005 ^ n13001 ;
  assign n13007 = n13002 & ~n13006 ;
  assign n13008 = n13007 ^ n11470 ;
  assign n13009 = n13008 ^ n11465 ;
  assign n13010 = ~n12116 & ~n12749 ;
  assign n13011 = n13010 ^ n12724 ;
  assign n13012 = n13011 ^ n13008 ;
  assign n13013 = n13009 & n13012 ;
  assign n13014 = n13013 ^ n11465 ;
  assign n13015 = n13014 ^ n10840 ;
  assign n13016 = n12751 ^ n12720 ;
  assign n13017 = ~n12113 & ~n13016 ;
  assign n13018 = n13017 ^ n12719 ;
  assign n13019 = n13018 ^ n13014 ;
  assign n13020 = ~n13015 & ~n13019 ;
  assign n13021 = n13020 ^ n10840 ;
  assign n13022 = n13021 ^ n11461 ;
  assign n13023 = n12109 & n12755 ;
  assign n13024 = n13023 ^ n12716 ;
  assign n13025 = n13024 ^ n13021 ;
  assign n13026 = ~n13022 & ~n13025 ;
  assign n13027 = n13026 ^ n11461 ;
  assign n13028 = n13027 ^ n12985 ;
  assign n13029 = n12986 & ~n13028 ;
  assign n13030 = n13029 ^ n10885 ;
  assign n13031 = n13030 ^ n12982 ;
  assign n13032 = n12983 & n13031 ;
  assign n13033 = n13032 ^ n10892 ;
  assign n13034 = n13033 ^ n12979 ;
  assign n13035 = n12980 & n13034 ;
  assign n13036 = n13035 ^ n11298 ;
  assign n13037 = n13036 ^ n12976 ;
  assign n13038 = n12977 & ~n13037 ;
  assign n13039 = n13038 ^ n10910 ;
  assign n13040 = n13039 ^ n10925 ;
  assign n13041 = ~n11643 & ~n12770 ;
  assign n13042 = n13041 ^ n12696 ;
  assign n13043 = n13042 ^ n13039 ;
  assign n13044 = ~n13040 & n13043 ;
  assign n13045 = n13044 ^ n10925 ;
  assign n13046 = n13045 ^ n10941 ;
  assign n13047 = ~n11638 & ~n12773 ;
  assign n13048 = n13047 ^ n12693 ;
  assign n13049 = n13048 ^ n13045 ;
  assign n13050 = n13046 & n13049 ;
  assign n13051 = n13050 ^ n10941 ;
  assign n13052 = n13051 ^ n12973 ;
  assign n13053 = n12974 & n13052 ;
  assign n13054 = n13053 ^ n10957 ;
  assign n13055 = n13054 ^ n12970 ;
  assign n13056 = n12971 & n13055 ;
  assign n13057 = n13056 ^ n10973 ;
  assign n13060 = n13059 ^ n13057 ;
  assign n13061 = n12966 ^ n10988 ;
  assign n13062 = n13061 ^ n12966 ;
  assign n13063 = n13062 ^ n13057 ;
  assign n13064 = n13060 & n13063 ;
  assign n13065 = n13064 ^ n13061 ;
  assign n13066 = n12967 & n13065 ;
  assign n13067 = n13066 ^ n11559 ;
  assign n13068 = n13067 ^ n11573 ;
  assign n13069 = n12227 & n12893 ;
  assign n13070 = n13069 ^ n12248 ;
  assign n13071 = n13070 ^ n13067 ;
  assign n13072 = ~n13068 & n13071 ;
  assign n13073 = n13072 ^ n11573 ;
  assign n13074 = n13073 ^ n12963 ;
  assign n13075 = n12964 & n13074 ;
  assign n13076 = n13075 ^ n11133 ;
  assign n13077 = n13076 ^ n12960 ;
  assign n13078 = ~n12961 & n13077 ;
  assign n13079 = n13078 ^ n11158 ;
  assign n13080 = n13079 ^ n11181 ;
  assign n12926 = n12433 ^ x7 ;
  assign n12923 = n12921 ^ n12281 ;
  assign n12924 = n12922 & n12923 ;
  assign n12810 = n12281 ^ n12276 ;
  assign n12925 = n12924 ^ n12810 ;
  assign n13081 = n12926 ^ n12925 ;
  assign n13082 = n13081 ^ n12276 ;
  assign n13083 = ~n11614 & n13082 ;
  assign n13084 = n13083 ^ n12276 ;
  assign n13085 = n13084 ^ n13079 ;
  assign n13086 = ~n13080 & n13085 ;
  assign n13087 = n13086 ^ n11181 ;
  assign n13088 = n13087 ^ n11204 ;
  assign n12927 = n12926 ^ n12276 ;
  assign n12928 = n12925 & n12927 ;
  assign n12809 = n12276 ^ n12271 ;
  assign n12929 = n12928 ^ n12809 ;
  assign n13089 = n12929 ^ n12613 ;
  assign n13090 = n13089 ^ n12271 ;
  assign n13091 = ~n11609 & n13090 ;
  assign n13092 = n13091 ^ n12271 ;
  assign n13093 = n13092 ^ n13087 ;
  assign n13094 = ~n13088 & ~n13093 ;
  assign n13095 = n13094 ^ n11204 ;
  assign n13096 = n13095 ^ n11227 ;
  assign n12935 = n12614 ^ n12613 ;
  assign n12931 = n12271 ^ n12266 ;
  assign n12930 = n12613 ^ n12266 ;
  assign n12932 = n12931 ^ n12930 ;
  assign n12933 = ~n12929 & n12932 ;
  assign n12934 = n12933 ^ n12930 ;
  assign n13097 = n12935 ^ n12934 ;
  assign n13098 = n13097 ^ n12266 ;
  assign n13099 = ~n11604 & n13098 ;
  assign n13100 = n13099 ^ n12266 ;
  assign n13101 = n13100 ^ n13095 ;
  assign n13102 = ~n13096 & n13101 ;
  assign n13103 = n13102 ^ n11227 ;
  assign n12940 = n12616 ^ n12615 ;
  assign n12938 = n12420 ^ n12266 ;
  assign n12936 = n12935 ^ n12266 ;
  assign n12937 = n12934 & n12936 ;
  assign n12939 = n12938 ^ n12937 ;
  assign n12955 = n12940 ^ n12939 ;
  assign n12956 = n12955 ^ n12420 ;
  assign n12957 = ~n11768 & n12956 ;
  assign n12958 = n12957 ^ n12420 ;
  assign n13104 = n13103 ^ n12958 ;
  assign n12941 = n12940 ^ n12420 ;
  assign n12942 = n12939 & n12941 ;
  assign n12943 = n12942 ^ n12420 ;
  assign n12808 = n12618 ^ n12617 ;
  assign n12944 = n12943 ^ n12808 ;
  assign n13105 = ~n11779 & n12944 ;
  assign n12945 = n12579 ^ n11779 ;
  assign n12946 = n12945 ^ n12582 ;
  assign n13106 = n13105 ^ n12946 ;
  assign n13107 = n13106 ^ n11242 ;
  assign n13108 = n13107 ^ n12958 ;
  assign n13109 = n13108 ^ n13106 ;
  assign n13110 = ~n13104 & ~n13109 ;
  assign n13111 = n13110 ^ n13107 ;
  assign n12950 = n12620 ^ n12619 ;
  assign n12947 = n12946 ^ n12808 ;
  assign n12948 = n12944 & ~n12947 ;
  assign n12949 = n12948 ^ n12943 ;
  assign n12951 = n12950 ^ n12949 ;
  assign n12952 = ~n12664 & ~n12951 ;
  assign n12953 = n12952 ^ n12601 ;
  assign n13113 = n12953 ^ n11775 ;
  assign n13112 = n13106 ^ n12953 ;
  assign n13114 = n13113 ^ n13112 ;
  assign n13115 = n13111 & n13114 ;
  assign n13116 = n13115 ^ n13113 ;
  assign n13131 = n13116 ^ n11331 ;
  assign n13132 = n13131 ^ x190 ;
  assign n13134 = n13103 ^ n11242 ;
  assign n13135 = n13134 ^ n12958 ;
  assign n13136 = n13135 ^ x176 ;
  assign n13138 = n13057 ^ n10988 ;
  assign n13139 = n13138 ^ n13059 ;
  assign n13140 = n13139 ^ x168 ;
  assign n13207 = n13042 ^ n13040 ;
  assign n13141 = n13036 ^ n10910 ;
  assign n13142 = n13141 ^ n12976 ;
  assign n13143 = n13142 ^ x173 ;
  assign n13145 = n12991 ^ n11475 ;
  assign n13146 = x167 & ~n13145 ;
  assign n13144 = n12996 ^ n11477 ;
  assign n13147 = n13146 ^ n13144 ;
  assign n13148 = n12998 ^ n11472 ;
  assign n13149 = n13148 ^ n12988 ;
  assign n13150 = n13149 ^ x166 ;
  assign n13151 = n13150 ^ n13146 ;
  assign n13152 = n13151 ^ n13149 ;
  assign n13153 = ~n13147 & n13152 ;
  assign n13154 = n13153 ^ n13150 ;
  assign n13155 = n13005 ^ n13002 ;
  assign n13157 = n13155 ^ x165 ;
  assign n13156 = n13155 ^ n13149 ;
  assign n13158 = n13157 ^ n13156 ;
  assign n13159 = ~n13154 & n13158 ;
  assign n13160 = n13159 ^ n13157 ;
  assign n13161 = n13011 ^ n13009 ;
  assign n13163 = n13161 ^ x164 ;
  assign n13162 = n13161 ^ n13155 ;
  assign n13164 = n13163 ^ n13162 ;
  assign n13165 = ~n13160 & n13164 ;
  assign n13166 = n13165 ^ n13163 ;
  assign n13167 = n13018 ^ n13015 ;
  assign n13169 = n13167 ^ x163 ;
  assign n13168 = n13167 ^ n13161 ;
  assign n13170 = n13169 ^ n13168 ;
  assign n13171 = n13166 & ~n13170 ;
  assign n13172 = n13171 ^ n13169 ;
  assign n13173 = n13024 ^ n13022 ;
  assign n13175 = n13173 ^ x162 ;
  assign n13174 = n13173 ^ n13167 ;
  assign n13176 = n13175 ^ n13174 ;
  assign n13177 = n13172 & ~n13176 ;
  assign n13178 = n13177 ^ n13175 ;
  assign n13179 = n13027 ^ n10885 ;
  assign n13180 = n13179 ^ n12985 ;
  assign n13182 = n13180 ^ x161 ;
  assign n13181 = n13180 ^ n13173 ;
  assign n13183 = n13182 ^ n13181 ;
  assign n13184 = ~n13178 & n13183 ;
  assign n13185 = n13184 ^ n13182 ;
  assign n13186 = n13030 ^ n10892 ;
  assign n13187 = n13186 ^ n12982 ;
  assign n13189 = n13187 ^ x160 ;
  assign n13188 = n13187 ^ n13180 ;
  assign n13190 = n13189 ^ n13188 ;
  assign n13191 = ~n13185 & n13190 ;
  assign n13192 = n13191 ^ n13189 ;
  assign n13193 = n13033 ^ n11298 ;
  assign n13194 = n13193 ^ n12979 ;
  assign n13196 = n13194 ^ x175 ;
  assign n13195 = n13194 ^ n13187 ;
  assign n13197 = n13196 ^ n13195 ;
  assign n13198 = ~n13192 & n13197 ;
  assign n13199 = n13198 ^ n13196 ;
  assign n13201 = n13142 ^ x174 ;
  assign n13200 = n13194 ^ n13142 ;
  assign n13202 = n13201 ^ n13200 ;
  assign n13203 = n13199 & ~n13202 ;
  assign n13204 = n13203 ^ n13201 ;
  assign n13205 = n13143 & ~n13204 ;
  assign n13206 = n13205 ^ x173 ;
  assign n13208 = n13207 ^ n13206 ;
  assign n13209 = n13048 ^ n13046 ;
  assign n13210 = n13209 ^ x172 ;
  assign n13211 = n13210 ^ n13206 ;
  assign n13212 = n13211 ^ n13209 ;
  assign n13213 = ~n13208 & n13212 ;
  assign n13214 = n13213 ^ n13210 ;
  assign n13215 = n13051 ^ n10957 ;
  assign n13216 = n13215 ^ n12973 ;
  assign n13218 = n13216 ^ x171 ;
  assign n13217 = n13216 ^ n13209 ;
  assign n13219 = n13218 ^ n13217 ;
  assign n13220 = ~n13214 & n13219 ;
  assign n13221 = n13220 ^ n13218 ;
  assign n13222 = n13054 ^ n10973 ;
  assign n13223 = n13222 ^ n12970 ;
  assign n13225 = n13223 ^ x170 ;
  assign n13224 = n13223 ^ n13216 ;
  assign n13226 = n13225 ^ n13224 ;
  assign n13227 = n13221 & ~n13226 ;
  assign n13228 = n13227 ^ n13225 ;
  assign n13230 = n13139 ^ x169 ;
  assign n13229 = n13223 ^ n13139 ;
  assign n13231 = n13230 ^ n13229 ;
  assign n13232 = ~n13228 & n13231 ;
  assign n13233 = n13232 ^ n13230 ;
  assign n13234 = n13140 & ~n13233 ;
  assign n13235 = n13234 ^ x168 ;
  assign n13137 = n13065 ^ n11559 ;
  assign n13236 = n13235 ^ n13137 ;
  assign n13237 = n13070 ^ n13068 ;
  assign n13238 = n13237 ^ x183 ;
  assign n13239 = n13238 ^ n13137 ;
  assign n13240 = n13239 ^ n13237 ;
  assign n13241 = n13236 & ~n13240 ;
  assign n13242 = n13241 ^ n13238 ;
  assign n13243 = n13073 ^ n11133 ;
  assign n13244 = n13243 ^ n12963 ;
  assign n13246 = n13244 ^ x182 ;
  assign n13245 = n13244 ^ n13237 ;
  assign n13247 = n13246 ^ n13245 ;
  assign n13248 = ~n13242 & n13247 ;
  assign n13249 = n13248 ^ n13246 ;
  assign n13250 = n13076 ^ n11158 ;
  assign n13251 = n13250 ^ n12960 ;
  assign n13253 = n13251 ^ x181 ;
  assign n13252 = n13251 ^ n13244 ;
  assign n13254 = n13253 ^ n13252 ;
  assign n13255 = n13249 & ~n13254 ;
  assign n13256 = n13255 ^ n13253 ;
  assign n13257 = n13084 ^ n13080 ;
  assign n13259 = n13257 ^ x180 ;
  assign n13258 = n13257 ^ n13251 ;
  assign n13260 = n13259 ^ n13258 ;
  assign n13261 = n13256 & ~n13260 ;
  assign n13262 = n13261 ^ n13259 ;
  assign n13263 = n13092 ^ n13088 ;
  assign n13265 = n13263 ^ x179 ;
  assign n13264 = n13263 ^ n13257 ;
  assign n13266 = n13265 ^ n13264 ;
  assign n13267 = ~n13262 & n13266 ;
  assign n13268 = n13267 ^ n13265 ;
  assign n13269 = n13100 ^ n13096 ;
  assign n13271 = n13269 ^ x178 ;
  assign n13270 = n13269 ^ n13263 ;
  assign n13272 = n13271 ^ n13270 ;
  assign n13273 = ~n13268 & n13272 ;
  assign n13274 = n13273 ^ n13271 ;
  assign n13276 = n13135 ^ x177 ;
  assign n13275 = n13269 ^ n13135 ;
  assign n13277 = n13276 ^ n13275 ;
  assign n13278 = ~n13274 & n13277 ;
  assign n13279 = n13278 ^ n13276 ;
  assign n13280 = n13136 & ~n13279 ;
  assign n13281 = n13280 ^ x176 ;
  assign n13133 = n13111 ^ n11775 ;
  assign n13282 = n13281 ^ n13133 ;
  assign n13283 = n13131 ^ x191 ;
  assign n13284 = n13283 ^ n13131 ;
  assign n13285 = n13284 ^ n13133 ;
  assign n13286 = ~n13282 & n13285 ;
  assign n13287 = n13286 ^ n13283 ;
  assign n13288 = ~n13132 & n13287 ;
  assign n13289 = n13288 ^ x190 ;
  assign n13120 = n12664 ^ n12601 ;
  assign n13121 = n13120 ^ n12949 ;
  assign n13122 = n12622 ^ n12621 ;
  assign n13123 = n13122 ^ n12950 ;
  assign n13124 = n13123 ^ n13122 ;
  assign n13125 = n13124 ^ n12949 ;
  assign n13126 = ~n13121 & n13125 ;
  assign n13127 = n13126 ^ n13123 ;
  assign n13128 = n11966 & n13127 ;
  assign n13129 = n13128 ^ n12670 ;
  assign n12954 = n12953 ^ n11331 ;
  assign n13117 = n12954 & n13116 ;
  assign n13118 = n13117 ^ n11331 ;
  assign n13119 = n13118 ^ n11959 ;
  assign n13130 = n13129 ^ n13119 ;
  assign n13290 = n13289 ^ n13130 ;
  assign n13301 = n12624 ^ n12623 ;
  assign n13297 = n12791 ^ n12670 ;
  assign n13296 = n13122 ^ n12791 ;
  assign n13298 = n13297 ^ n13296 ;
  assign n13299 = ~n13127 & n13298 ;
  assign n13300 = n13299 ^ n13297 ;
  assign n13302 = n13301 ^ n13300 ;
  assign n13303 = n13302 ^ n12791 ;
  assign n13304 = n12784 & n13303 ;
  assign n13305 = n13304 ^ n12791 ;
  assign n13291 = n13129 ^ n13118 ;
  assign n13292 = n13129 ^ n11959 ;
  assign n13293 = n13291 & ~n13292 ;
  assign n13294 = n13293 ^ n11959 ;
  assign n13295 = n13294 ^ n11370 ;
  assign n13306 = n13305 ^ n13295 ;
  assign n13307 = n13306 ^ x189 ;
  assign n13308 = n13307 ^ n13289 ;
  assign n13309 = n13308 ^ n13306 ;
  assign n13310 = n13290 & n13309 ;
  assign n13311 = n13310 ^ n13307 ;
  assign n13432 = n13311 ^ x188 ;
  assign n13376 = n13214 ^ x171 ;
  assign n13377 = n13145 ^ x167 ;
  assign n13378 = n13147 ^ x166 ;
  assign n13379 = ~n13377 & n13378 ;
  assign n13380 = n13154 ^ x165 ;
  assign n13381 = ~n13379 & ~n13380 ;
  assign n13382 = n13160 ^ x164 ;
  assign n13383 = n13381 & ~n13382 ;
  assign n13384 = n13166 ^ x163 ;
  assign n13385 = n13383 & n13384 ;
  assign n13386 = n13172 ^ x162 ;
  assign n13387 = ~n13385 & ~n13386 ;
  assign n13388 = n13178 ^ x161 ;
  assign n13389 = ~n13387 & ~n13388 ;
  assign n13390 = n13185 ^ x160 ;
  assign n13391 = ~n13389 & n13390 ;
  assign n13392 = n13192 ^ x175 ;
  assign n13393 = n13391 & n13392 ;
  assign n13394 = n13199 ^ x174 ;
  assign n13395 = n13393 & ~n13394 ;
  assign n13396 = n13204 ^ x173 ;
  assign n13397 = n13395 & n13396 ;
  assign n13398 = n13206 ^ x172 ;
  assign n13399 = n13398 ^ n13207 ;
  assign n13400 = n13397 & n13399 ;
  assign n13401 = ~n13376 & ~n13400 ;
  assign n13402 = n13221 ^ x170 ;
  assign n13403 = ~n13401 & ~n13402 ;
  assign n13404 = n13228 ^ x169 ;
  assign n13405 = n13403 & n13404 ;
  assign n13406 = n13233 ^ x168 ;
  assign n13407 = n13405 & n13406 ;
  assign n13408 = n13235 ^ x183 ;
  assign n13409 = n13408 ^ n13137 ;
  assign n13410 = ~n13407 & n13409 ;
  assign n13411 = n13242 ^ x182 ;
  assign n13412 = n13410 & ~n13411 ;
  assign n13413 = n13249 ^ x181 ;
  assign n13414 = n13412 & n13413 ;
  assign n13415 = n13256 ^ x180 ;
  assign n13416 = n13414 & n13415 ;
  assign n13417 = n13262 ^ x179 ;
  assign n13418 = ~n13416 & n13417 ;
  assign n13419 = n13268 ^ x178 ;
  assign n13420 = ~n13418 & ~n13419 ;
  assign n13421 = n13274 ^ x177 ;
  assign n13422 = ~n13420 & n13421 ;
  assign n13423 = n13279 ^ x176 ;
  assign n13424 = n13422 & n13423 ;
  assign n13425 = n13281 ^ x191 ;
  assign n13426 = n13425 ^ n13133 ;
  assign n13427 = n13424 & n13426 ;
  assign n13428 = n13287 ^ x190 ;
  assign n13429 = ~n13427 & n13428 ;
  assign n13430 = n13290 ^ x189 ;
  assign n13431 = n13429 & n13430 ;
  assign n13472 = n13432 ^ n13431 ;
  assign n13471 = n12735 ^ n12734 ;
  assign n14134 = n13472 ^ n13471 ;
  assign n13568 = n12735 & ~n13472 ;
  assign n13569 = n13568 ^ n12734 ;
  assign n13575 = n13569 ^ n12125 ;
  assign n13576 = x327 & ~n13575 ;
  assign n13322 = n12626 ^ n12625 ;
  assign n13318 = n12820 ^ n12791 ;
  assign n13317 = n13301 ^ n12820 ;
  assign n13319 = n13318 ^ n13317 ;
  assign n13320 = n13300 & n13319 ;
  assign n13321 = n13320 ^ n13318 ;
  assign n13323 = n13322 ^ n13321 ;
  assign n13324 = n13323 ^ n12820 ;
  assign n13325 = ~n12006 & n13324 ;
  assign n13326 = n13325 ^ n12820 ;
  assign n13312 = n13305 ^ n13294 ;
  assign n13313 = n13305 ^ n11370 ;
  assign n13314 = n13312 & ~n13313 ;
  assign n13315 = n13314 ^ n11370 ;
  assign n13316 = n13315 ^ n11391 ;
  assign n13327 = n13326 ^ n13316 ;
  assign n13329 = n13327 ^ x188 ;
  assign n13328 = n13327 ^ n13306 ;
  assign n13330 = n13329 ^ n13328 ;
  assign n13331 = n13311 & ~n13330 ;
  assign n13332 = n13331 ^ n13329 ;
  assign n13434 = n13332 ^ x187 ;
  assign n13433 = ~n13431 & ~n13432 ;
  assign n13476 = n13434 ^ n13433 ;
  assign n13473 = n13471 & n13472 ;
  assign n13477 = n13476 ^ n13473 ;
  assign n13572 = n12737 & n13477 ;
  assign n13474 = n12739 ^ n12738 ;
  assign n13573 = n13572 ^ n13474 ;
  assign n13570 = ~n12125 & n13569 ;
  assign n13571 = n13570 ^ n12128 ;
  assign n13574 = n13573 ^ n13571 ;
  assign n13577 = n13576 ^ n13574 ;
  assign n13475 = n13474 ^ n13473 ;
  assign n13478 = ~n13475 & ~n13477 ;
  assign n13479 = n13478 ^ n13474 ;
  assign n13343 = n12628 ^ n12627 ;
  assign n13339 = n12840 ^ n12820 ;
  assign n13338 = n13322 ^ n12840 ;
  assign n13340 = n13339 ^ n13338 ;
  assign n13341 = n13321 & n13340 ;
  assign n13342 = n13341 ^ n13339 ;
  assign n13344 = n13343 ^ n13342 ;
  assign n13345 = n13344 ^ n12840 ;
  assign n13346 = ~n12833 & ~n13345 ;
  assign n13347 = n13346 ^ n12840 ;
  assign n13333 = n13326 ^ n13315 ;
  assign n13334 = n13326 ^ n11391 ;
  assign n13335 = n13333 & ~n13334 ;
  assign n13336 = n13335 ^ n11391 ;
  assign n13337 = n13336 ^ n11408 ;
  assign n13348 = n13347 ^ n13337 ;
  assign n13350 = n13348 ^ x187 ;
  assign n13349 = n13348 ^ n13327 ;
  assign n13351 = n13350 ^ n13349 ;
  assign n13352 = n13332 & ~n13351 ;
  assign n13353 = n13352 ^ n13350 ;
  assign n13436 = n13353 ^ x186 ;
  assign n13435 = ~n13433 & n13434 ;
  assign n13469 = n13436 ^ n13435 ;
  assign n13582 = n13479 ^ n13469 ;
  assign n13583 = n12732 & n13582 ;
  assign n13467 = n12742 ^ n12732 ;
  assign n13468 = n13467 ^ n12730 ;
  assign n13584 = n13583 ^ n13468 ;
  assign n13578 = n13573 ^ n13570 ;
  assign n13579 = n13571 & n13578 ;
  assign n13580 = n13579 ^ n12128 ;
  assign n13581 = n13580 ^ n12123 ;
  assign n13585 = n13584 ^ n13581 ;
  assign n13586 = n13585 ^ x326 ;
  assign n13587 = n13586 ^ n13574 ;
  assign n13588 = n13587 ^ n13585 ;
  assign n13589 = n13577 & ~n13588 ;
  assign n13590 = n13589 ^ n13586 ;
  assign n13470 = n13469 ^ n13468 ;
  assign n13480 = n13479 ^ n13468 ;
  assign n13481 = ~n13470 & n13480 ;
  assign n13482 = n13481 ^ n13469 ;
  assign n13364 = n12630 ^ n12629 ;
  assign n13360 = n12867 ^ n12840 ;
  assign n13359 = n13343 ^ n12867 ;
  assign n13361 = n13360 ^ n13359 ;
  assign n13362 = ~n13342 & n13361 ;
  assign n13363 = n13362 ^ n13360 ;
  assign n13365 = n13364 ^ n13363 ;
  assign n13366 = n13365 ^ n12867 ;
  assign n13367 = n12176 & n13366 ;
  assign n13368 = n13367 ^ n12867 ;
  assign n13354 = n13347 ^ n13336 ;
  assign n13355 = n13347 ^ n11408 ;
  assign n13356 = ~n13354 & n13355 ;
  assign n13357 = n13356 ^ n11408 ;
  assign n13358 = n13357 ^ n11433 ;
  assign n13369 = n13368 ^ n13358 ;
  assign n13371 = n13369 ^ x186 ;
  assign n13370 = n13369 ^ n13348 ;
  assign n13372 = n13371 ^ n13370 ;
  assign n13373 = ~n13353 & n13372 ;
  assign n13374 = n13373 ^ n13371 ;
  assign n13463 = n13374 ^ x185 ;
  assign n13437 = ~n13435 & n13436 ;
  assign n13464 = n13463 ^ n13437 ;
  assign n13483 = n13482 ^ n13464 ;
  assign n13595 = n12727 & n13483 ;
  assign n13465 = n12746 ^ n12728 ;
  assign n13596 = n13595 ^ n13465 ;
  assign n13591 = n13584 ^ n13580 ;
  assign n13592 = ~n13581 & ~n13591 ;
  assign n13593 = n13592 ^ n12123 ;
  assign n13594 = n13593 ^ n12120 ;
  assign n13597 = n13596 ^ n13594 ;
  assign n13599 = n13597 ^ x325 ;
  assign n13598 = n13597 ^ n13585 ;
  assign n13600 = n13599 ^ n13598 ;
  assign n13601 = n13590 & ~n13600 ;
  assign n13602 = n13601 ^ n13599 ;
  assign n13466 = n13465 ^ n13464 ;
  assign n13484 = n13466 & ~n13483 ;
  assign n13485 = n13484 ^ n13465 ;
  assign n13453 = n13364 ^ n12867 ;
  assign n13454 = n13363 & ~n13453 ;
  assign n13450 = n12917 ^ n12631 ;
  assign n13451 = n13450 ^ n12632 ;
  assign n13452 = n13451 ^ n13364 ;
  assign n13455 = n13454 ^ n13452 ;
  assign n13456 = n13455 ^ n12917 ;
  assign n13457 = ~n12206 & n13456 ;
  assign n13447 = n12917 ^ n11509 ;
  assign n13446 = n11433 ^ x184 ;
  assign n13448 = n13447 ^ n13446 ;
  assign n13443 = n13368 ^ n13357 ;
  assign n13444 = n13368 ^ n11433 ;
  assign n13445 = n13443 & n13444 ;
  assign n13449 = n13448 ^ n13445 ;
  assign n13458 = n13457 ^ n13449 ;
  assign n13438 = n13437 ^ n13369 ;
  assign n13441 = ~n13374 & ~n13438 ;
  assign n13375 = n13374 ^ n13369 ;
  assign n13439 = n13438 ^ n13375 ;
  assign n13440 = x185 & ~n13439 ;
  assign n13442 = n13441 ^ n13440 ;
  assign n13459 = n13458 ^ n13442 ;
  assign n13486 = n13485 ^ n13459 ;
  assign n13607 = ~n12724 & n13486 ;
  assign n13460 = n12748 ^ n12724 ;
  assign n13461 = n13460 ^ n12722 ;
  assign n13608 = n13607 ^ n13461 ;
  assign n13603 = n13596 ^ n13593 ;
  assign n13604 = ~n13594 & ~n13603 ;
  assign n13605 = n13604 ^ n12120 ;
  assign n13606 = n13605 ^ n12116 ;
  assign n13609 = n13608 ^ n13606 ;
  assign n13611 = n13609 ^ x324 ;
  assign n13610 = n13609 ^ n13597 ;
  assign n13612 = n13611 ^ n13610 ;
  assign n13613 = ~n13602 & n13612 ;
  assign n13614 = n13613 ^ n13611 ;
  assign n13462 = n13461 ^ n13459 ;
  assign n13487 = ~n13462 & ~n13486 ;
  assign n13488 = n13487 ^ n13461 ;
  assign n13619 = n13488 ^ n13377 ;
  assign n13620 = n12719 & n13619 ;
  assign n13489 = n12752 ^ n12720 ;
  assign n13621 = n13620 ^ n13489 ;
  assign n13615 = n13608 ^ n13605 ;
  assign n13616 = ~n13606 & ~n13615 ;
  assign n13617 = n13616 ^ n12116 ;
  assign n13618 = n13617 ^ n12113 ;
  assign n13622 = n13621 ^ n13618 ;
  assign n13624 = n13622 ^ x323 ;
  assign n13623 = n13622 ^ n13609 ;
  assign n13625 = n13624 ^ n13623 ;
  assign n13626 = n13614 & ~n13625 ;
  assign n13627 = n13626 ^ n13624 ;
  assign n13628 = n13627 ^ x322 ;
  assign n13629 = n13590 ^ x325 ;
  assign n13630 = n13575 ^ x327 ;
  assign n13631 = n13576 ^ x326 ;
  assign n13632 = n13631 ^ n13574 ;
  assign n13633 = n13630 & n13632 ;
  assign n13634 = ~n13629 & ~n13633 ;
  assign n13635 = n13602 ^ x324 ;
  assign n13636 = n13634 & n13635 ;
  assign n13637 = n13614 ^ x323 ;
  assign n13638 = ~n13636 & n13637 ;
  assign n14055 = ~n13628 & ~n13638 ;
  assign n13858 = n13622 ^ x322 ;
  assign n13859 = n13627 & ~n13858 ;
  assign n13860 = n13859 ^ x322 ;
  assign n13701 = n13621 ^ n13617 ;
  assign n13702 = n13618 & ~n13701 ;
  assign n13703 = n13702 ^ n12113 ;
  assign n13705 = n13703 ^ n12109 ;
  assign n13498 = n13378 ^ n13377 ;
  assign n13490 = n13489 ^ n13488 ;
  assign n13491 = n12754 ^ n12716 ;
  assign n13492 = n13491 ^ n12714 ;
  assign n13493 = n13492 ^ n13377 ;
  assign n13494 = n13493 ^ n13492 ;
  assign n13495 = n13494 ^ n13488 ;
  assign n13496 = n13490 & n13495 ;
  assign n13497 = n13496 ^ n13493 ;
  assign n13697 = n13498 ^ n13497 ;
  assign n13698 = n13697 ^ n13492 ;
  assign n13699 = ~n12716 & ~n13698 ;
  assign n13700 = n13699 ^ n13492 ;
  assign n13857 = n13705 ^ n13700 ;
  assign n13861 = n13860 ^ n13857 ;
  assign n14056 = n13861 ^ x321 ;
  assign n14057 = ~n14055 & ~n14056 ;
  assign n13704 = n13703 ^ n13700 ;
  assign n13706 = ~n13704 & ~n13705 ;
  assign n13707 = n13706 ^ n12109 ;
  assign n13709 = n13707 ^ n12105 ;
  assign n13506 = n13380 ^ n13379 ;
  assign n13499 = n12757 ^ n12712 ;
  assign n13500 = n13499 ^ n12710 ;
  assign n13502 = n13500 ^ n13492 ;
  assign n13501 = n13500 ^ n13498 ;
  assign n13503 = n13502 ^ n13501 ;
  assign n13504 = ~n13497 & n13503 ;
  assign n13505 = n13504 ^ n13502 ;
  assign n13693 = n13506 ^ n13505 ;
  assign n13694 = n13693 ^ n13500 ;
  assign n13695 = n12712 & n13694 ;
  assign n13696 = n13695 ^ n13500 ;
  assign n13862 = n13709 ^ n13696 ;
  assign n13863 = n13862 ^ x321 ;
  assign n13864 = n13863 ^ n13860 ;
  assign n13865 = n13864 ^ n13862 ;
  assign n13866 = ~n13861 & n13865 ;
  assign n13867 = n13866 ^ n13863 ;
  assign n14058 = n13867 ^ x320 ;
  assign n14059 = ~n14057 & ~n14058 ;
  assign n13708 = n13707 ^ n13696 ;
  assign n13710 = n13708 & n13709 ;
  assign n13711 = n13710 ^ n12105 ;
  assign n13868 = n13711 ^ n12101 ;
  assign n13514 = n13382 ^ n13381 ;
  assign n13507 = n12760 ^ n12708 ;
  assign n13508 = n13507 ^ n12706 ;
  assign n13510 = n13508 ^ n13500 ;
  assign n13509 = n13508 ^ n13506 ;
  assign n13511 = n13510 ^ n13509 ;
  assign n13512 = n13505 & n13511 ;
  assign n13513 = n13512 ^ n13510 ;
  assign n13688 = n13514 ^ n13513 ;
  assign n13689 = n13688 ^ n13508 ;
  assign n13690 = ~n12708 & ~n13689 ;
  assign n13691 = n13690 ^ n13508 ;
  assign n13869 = n13868 ^ n13691 ;
  assign n13871 = n13869 ^ x320 ;
  assign n13870 = n13869 ^ n13862 ;
  assign n13872 = n13871 ^ n13870 ;
  assign n13873 = n13867 & ~n13872 ;
  assign n13874 = n13873 ^ n13871 ;
  assign n14060 = n13874 ^ x335 ;
  assign n14061 = n14059 & n14060 ;
  assign n13692 = n13691 ^ n12101 ;
  assign n13712 = n13711 ^ n13691 ;
  assign n13713 = n13692 & ~n13712 ;
  assign n13714 = n13713 ^ n12101 ;
  assign n13875 = n13714 ^ n11705 ;
  assign n13522 = n13384 ^ n13383 ;
  assign n13515 = n12763 ^ n12704 ;
  assign n13516 = n13515 ^ n12702 ;
  assign n13518 = n13516 ^ n13508 ;
  assign n13517 = n13516 ^ n13514 ;
  assign n13519 = n13518 ^ n13517 ;
  assign n13520 = ~n13513 & n13519 ;
  assign n13521 = n13520 ^ n13518 ;
  assign n13683 = n13522 ^ n13521 ;
  assign n13684 = n13683 ^ n13516 ;
  assign n13685 = n12704 & ~n13684 ;
  assign n13686 = n13685 ^ n13516 ;
  assign n13876 = n13875 ^ n13686 ;
  assign n13878 = n13876 ^ x335 ;
  assign n13877 = n13876 ^ n13869 ;
  assign n13879 = n13878 ^ n13877 ;
  assign n13880 = ~n13874 & n13879 ;
  assign n13881 = n13880 ^ n13878 ;
  assign n14062 = n13881 ^ x334 ;
  assign n14063 = n14061 & ~n14062 ;
  assign n13687 = n13686 ^ n11705 ;
  assign n13715 = n13714 ^ n13686 ;
  assign n13716 = ~n13687 & ~n13715 ;
  assign n13717 = n13716 ^ n11705 ;
  assign n13882 = n13717 ^ n11648 ;
  assign n13530 = n13386 ^ n13385 ;
  assign n13523 = n12766 ^ n12700 ;
  assign n13524 = n13523 ^ n12698 ;
  assign n13526 = n13524 ^ n13516 ;
  assign n13525 = n13524 ^ n13522 ;
  assign n13527 = n13526 ^ n13525 ;
  assign n13528 = n13521 & ~n13527 ;
  assign n13529 = n13528 ^ n13526 ;
  assign n13646 = n13530 ^ n13529 ;
  assign n13679 = n13646 ^ n13524 ;
  assign n13680 = n12700 & n13679 ;
  assign n13681 = n13680 ^ n13524 ;
  assign n13883 = n13882 ^ n13681 ;
  assign n13885 = n13883 ^ x334 ;
  assign n13884 = n13883 ^ n13876 ;
  assign n13886 = n13885 ^ n13884 ;
  assign n13887 = n13881 & ~n13886 ;
  assign n13888 = n13887 ^ n13885 ;
  assign n14064 = n13888 ^ x333 ;
  assign n14065 = ~n14063 & ~n14064 ;
  assign n13682 = n13681 ^ n11648 ;
  assign n13718 = n13717 ^ n13681 ;
  assign n13719 = ~n13682 & ~n13718 ;
  assign n13720 = n13719 ^ n11648 ;
  assign n13889 = n13720 ^ n11643 ;
  assign n13538 = n13388 ^ n13387 ;
  assign n13531 = n12769 ^ n12696 ;
  assign n13532 = n13531 ^ n12695 ;
  assign n13534 = n13532 ^ n13524 ;
  assign n13533 = n13532 ^ n13530 ;
  assign n13535 = n13534 ^ n13533 ;
  assign n13536 = ~n13529 & ~n13535 ;
  assign n13537 = n13536 ^ n13534 ;
  assign n13647 = n13538 ^ n13537 ;
  assign n13675 = n13647 ^ n13532 ;
  assign n13676 = ~n12696 & n13675 ;
  assign n13677 = n13676 ^ n13532 ;
  assign n13890 = n13889 ^ n13677 ;
  assign n13892 = n13890 ^ x333 ;
  assign n13891 = n13890 ^ n13883 ;
  assign n13893 = n13892 ^ n13891 ;
  assign n13894 = ~n13888 & n13893 ;
  assign n13895 = n13894 ^ n13892 ;
  assign n14066 = n13895 ^ x332 ;
  assign n14067 = ~n14065 & ~n14066 ;
  assign n13547 = n13390 ^ n13389 ;
  assign n13539 = n12773 ^ n12693 ;
  assign n13541 = n13539 ^ n13532 ;
  assign n13540 = n13539 ^ n13538 ;
  assign n13542 = n13541 ^ n13540 ;
  assign n13543 = ~n13537 & ~n13542 ;
  assign n13544 = n13543 ^ n13541 ;
  assign n13641 = n13547 ^ n13544 ;
  assign n13725 = n13641 ^ n12773 ;
  assign n13726 = ~n12693 & ~n13725 ;
  assign n13727 = n13726 ^ n13641 ;
  assign n13678 = n13677 ^ n11643 ;
  assign n13721 = n13720 ^ n13677 ;
  assign n13722 = ~n13678 & ~n13721 ;
  assign n13723 = n13722 ^ n11643 ;
  assign n13724 = n13723 ^ n11638 ;
  assign n13896 = n13727 ^ n13724 ;
  assign n13898 = n13896 ^ x332 ;
  assign n13897 = n13896 ^ n13890 ;
  assign n13899 = n13898 ^ n13897 ;
  assign n13900 = n13895 & ~n13899 ;
  assign n13901 = n13900 ^ n13898 ;
  assign n14068 = n13901 ^ x331 ;
  assign n14069 = ~n14067 & ~n14068 ;
  assign n13728 = n13727 ^ n13723 ;
  assign n13729 = n13724 & n13728 ;
  assign n13730 = n13729 ^ n11638 ;
  assign n13902 = n13730 ^ n11633 ;
  assign n13553 = n13392 ^ n13391 ;
  assign n13545 = n12775 ^ n12689 ;
  assign n13546 = n13545 ^ n12688 ;
  assign n13549 = n13546 ^ n13539 ;
  assign n13548 = n13547 ^ n13546 ;
  assign n13550 = n13549 ^ n13548 ;
  assign n13551 = ~n13544 & n13550 ;
  assign n13552 = n13551 ^ n13549 ;
  assign n13642 = n13553 ^ n13552 ;
  assign n13671 = n13642 ^ n13546 ;
  assign n13672 = n12689 & ~n13671 ;
  assign n13673 = n13672 ^ n13546 ;
  assign n13903 = n13902 ^ n13673 ;
  assign n13905 = n13903 ^ x331 ;
  assign n13904 = n13903 ^ n13896 ;
  assign n13906 = n13905 ^ n13904 ;
  assign n13907 = ~n13901 & n13906 ;
  assign n13908 = n13907 ^ n13905 ;
  assign n14070 = n13908 ^ x330 ;
  assign n14071 = ~n14069 & n14070 ;
  assign n13674 = n13673 ^ n11633 ;
  assign n13731 = n13730 ^ n13673 ;
  assign n13732 = ~n13674 & ~n13731 ;
  assign n13733 = n13732 ^ n11633 ;
  assign n13909 = n13733 ^ n11556 ;
  assign n13556 = n13394 ^ n13393 ;
  assign n13557 = n13556 ^ n13546 ;
  assign n13554 = n13553 ^ n13546 ;
  assign n13555 = n13552 & ~n13554 ;
  assign n13558 = n13557 ^ n13555 ;
  assign n13668 = ~n12219 & n13558 ;
  assign n13559 = n12779 ^ n12686 ;
  assign n13669 = n13668 ^ n13559 ;
  assign n13910 = n13909 ^ n13669 ;
  assign n13912 = n13910 ^ x330 ;
  assign n13911 = n13910 ^ n13903 ;
  assign n13913 = n13912 ^ n13911 ;
  assign n13914 = ~n13908 & n13913 ;
  assign n13915 = n13914 ^ n13912 ;
  assign n14072 = n13915 ^ x329 ;
  assign n14073 = n14071 & ~n14072 ;
  assign n13670 = n13669 ^ n11556 ;
  assign n13734 = n13733 ^ n13669 ;
  assign n13735 = ~n13670 & ~n13734 ;
  assign n13736 = n13735 ^ n11556 ;
  assign n13854 = n13736 ^ n12231 ;
  assign n13565 = n13396 ^ n13395 ;
  assign n12782 = n12781 ^ n12384 ;
  assign n12807 = n12806 ^ n12782 ;
  assign n13563 = n13559 ^ n12807 ;
  assign n13561 = n13559 ^ n13556 ;
  assign n13562 = ~n13558 & ~n13561 ;
  assign n13564 = n13563 ^ n13562 ;
  assign n13566 = n13565 ^ n13564 ;
  assign n13737 = n13566 ^ n12807 ;
  assign n13738 = n12384 & n13737 ;
  assign n13739 = n13738 ^ n12807 ;
  assign n13855 = n13854 ^ n13739 ;
  assign n13917 = n13855 ^ x329 ;
  assign n13916 = n13910 ^ n13855 ;
  assign n13918 = n13917 ^ n13916 ;
  assign n13919 = n13915 & ~n13918 ;
  assign n13920 = n13919 ^ n13917 ;
  assign n14074 = n13920 ^ x328 ;
  assign n14075 = n14073 & ~n14074 ;
  assign n13856 = n13855 ^ x328 ;
  assign n13921 = ~n13856 & n13920 ;
  assign n13922 = n13921 ^ x328 ;
  assign n14076 = n13922 ^ x343 ;
  assign n13740 = n13739 ^ n13736 ;
  assign n13656 = n13399 ^ n13397 ;
  assign n13653 = n13565 ^ n12807 ;
  assign n13654 = ~n13564 & n13653 ;
  assign n13655 = n13654 ^ n13565 ;
  assign n13657 = n13656 ^ n13655 ;
  assign n13741 = ~n12884 & n13657 ;
  assign n13659 = n12889 ^ n12885 ;
  assign n13742 = n13741 ^ n13659 ;
  assign n13743 = n13742 ^ n12231 ;
  assign n13744 = n13743 ^ n13736 ;
  assign n13745 = n13744 ^ n13742 ;
  assign n13746 = n13740 & ~n13745 ;
  assign n13747 = n13746 ^ n13743 ;
  assign n13923 = n13747 ^ n12244 ;
  assign n14077 = n14076 ^ n13923 ;
  assign n14078 = n14075 & n14077 ;
  assign n13924 = n13923 ^ n13922 ;
  assign n13662 = n13659 ^ n13655 ;
  assign n13663 = ~n13657 & ~n13662 ;
  assign n13658 = n13400 ^ n13376 ;
  assign n13660 = n13659 ^ n13658 ;
  assign n13664 = n13663 ^ n13660 ;
  assign n13665 = ~n12881 & n13664 ;
  assign n13651 = n12892 ^ n12881 ;
  assign n13652 = n13651 ^ n12880 ;
  assign n13666 = n13665 ^ n13652 ;
  assign n13749 = n13666 ^ n12244 ;
  assign n13748 = n13742 ^ n13666 ;
  assign n13750 = n13749 ^ n13748 ;
  assign n13751 = n13747 & n13750 ;
  assign n13752 = n13751 ^ n13749 ;
  assign n13852 = n13752 ^ n12227 ;
  assign n13925 = n13852 ^ x343 ;
  assign n13926 = n13925 ^ n13852 ;
  assign n13927 = n13926 ^ n13922 ;
  assign n13928 = ~n13924 & n13927 ;
  assign n13929 = n13928 ^ n13925 ;
  assign n14079 = n13929 ^ x342 ;
  assign n14080 = n14078 & ~n14079 ;
  assign n13853 = n13852 ^ x342 ;
  assign n13930 = ~n13853 & n13929 ;
  assign n13931 = n13930 ^ x342 ;
  assign n14081 = n13931 ^ x341 ;
  assign n13758 = n13402 ^ n13401 ;
  assign n13760 = n13758 ^ n13658 ;
  assign n13759 = n13758 ^ n13652 ;
  assign n13761 = n13760 ^ n13759 ;
  assign n13762 = n13664 & ~n13761 ;
  assign n13763 = n13762 ^ n13760 ;
  assign n13764 = n12286 & ~n13763 ;
  assign n13756 = n12895 ^ n12286 ;
  assign n13757 = n13756 ^ n12878 ;
  assign n13765 = n13764 ^ n13757 ;
  assign n13667 = n13666 ^ n12227 ;
  assign n13753 = n13667 & n13752 ;
  assign n13754 = n13753 ^ n12227 ;
  assign n13755 = n13754 ^ n11624 ;
  assign n13932 = n13765 ^ n13755 ;
  assign n14082 = n14081 ^ n13932 ;
  assign n14083 = ~n14080 & n14082 ;
  assign n13933 = n13932 ^ n13931 ;
  assign n13777 = n13404 ^ n13403 ;
  assign n13770 = n12898 ^ n12281 ;
  assign n13771 = n13770 ^ n12921 ;
  assign n13773 = n13771 ^ n13757 ;
  assign n13772 = n13771 ^ n13758 ;
  assign n13774 = n13773 ^ n13772 ;
  assign n13775 = ~n13763 & n13774 ;
  assign n13776 = n13775 ^ n13772 ;
  assign n13778 = n13777 ^ n13776 ;
  assign n13779 = n13778 ^ n13771 ;
  assign n13780 = ~n12281 & n13779 ;
  assign n13781 = n13780 ^ n13771 ;
  assign n13766 = n13765 ^ n13754 ;
  assign n13767 = ~n13755 & ~n13766 ;
  assign n13768 = n13767 ^ n11624 ;
  assign n13769 = n13768 ^ n11619 ;
  assign n13934 = n13781 ^ n13769 ;
  assign n13935 = n13934 ^ x341 ;
  assign n13936 = n13935 ^ n13931 ;
  assign n13937 = n13936 ^ n13934 ;
  assign n13938 = n13933 & n13937 ;
  assign n13939 = n13938 ^ n13935 ;
  assign n14084 = n13939 ^ x340 ;
  assign n14085 = ~n14083 & ~n14084 ;
  assign n13786 = n13406 ^ n13405 ;
  assign n13788 = n13786 ^ n13771 ;
  assign n13787 = n13786 ^ n13777 ;
  assign n13789 = n13788 ^ n13787 ;
  assign n13790 = n13776 & n13789 ;
  assign n13791 = n13790 ^ n13788 ;
  assign n13792 = ~n12276 & n13791 ;
  assign n13793 = n13792 ^ n13081 ;
  assign n13782 = n13781 ^ n13768 ;
  assign n13783 = ~n13769 & n13782 ;
  assign n13784 = n13783 ^ n11619 ;
  assign n13785 = n13784 ^ n11614 ;
  assign n13940 = n13793 ^ n13785 ;
  assign n13942 = n13940 ^ x340 ;
  assign n13941 = n13940 ^ n13934 ;
  assign n13943 = n13942 ^ n13941 ;
  assign n13944 = n13939 & ~n13943 ;
  assign n13945 = n13944 ^ n13942 ;
  assign n14086 = n13945 ^ x339 ;
  assign n14087 = n14085 & n14086 ;
  assign n13803 = n13409 ^ n13407 ;
  assign n13799 = n13089 ^ n13081 ;
  assign n13798 = n13786 ^ n13089 ;
  assign n13800 = n13799 ^ n13798 ;
  assign n13801 = ~n13791 & ~n13800 ;
  assign n13802 = n13801 ^ n13799 ;
  assign n13804 = n13803 ^ n13802 ;
  assign n13805 = n13804 ^ n13089 ;
  assign n13806 = ~n12271 & ~n13805 ;
  assign n13807 = n13806 ^ n13089 ;
  assign n13794 = n13793 ^ n13784 ;
  assign n13795 = ~n13785 & n13794 ;
  assign n13796 = n13795 ^ n11614 ;
  assign n13797 = n13796 ^ n11609 ;
  assign n13946 = n13807 ^ n13797 ;
  assign n13948 = n13946 ^ x339 ;
  assign n13947 = n13946 ^ n13940 ;
  assign n13949 = n13948 ^ n13947 ;
  assign n13950 = ~n13945 & n13949 ;
  assign n13951 = n13950 ^ n13948 ;
  assign n14088 = n13951 ^ x338 ;
  assign n14089 = n14087 & ~n14088 ;
  assign n13817 = n13411 ^ n13410 ;
  assign n13813 = n13097 ^ n13089 ;
  assign n13812 = n13803 ^ n13097 ;
  assign n13814 = n13813 ^ n13812 ;
  assign n13815 = n13802 & ~n13814 ;
  assign n13816 = n13815 ^ n13813 ;
  assign n13818 = n13817 ^ n13816 ;
  assign n13819 = n13818 ^ n13097 ;
  assign n13820 = ~n12266 & ~n13819 ;
  assign n13821 = n13820 ^ n13097 ;
  assign n13808 = n13807 ^ n13796 ;
  assign n13809 = n13797 & ~n13808 ;
  assign n13810 = n13809 ^ n11609 ;
  assign n13811 = n13810 ^ n11604 ;
  assign n13952 = n13821 ^ n13811 ;
  assign n13954 = n13952 ^ x338 ;
  assign n13953 = n13952 ^ n13946 ;
  assign n13955 = n13954 ^ n13953 ;
  assign n13956 = n13951 & ~n13955 ;
  assign n13957 = n13956 ^ n13954 ;
  assign n14090 = n13957 ^ x337 ;
  assign n14091 = ~n14089 & n14090 ;
  assign n13822 = n13821 ^ n13810 ;
  assign n13823 = n13811 & ~n13822 ;
  assign n13824 = n13823 ^ n11604 ;
  assign n13849 = n13824 ^ n11768 ;
  assign n13830 = n13413 ^ n13412 ;
  assign n13826 = n13097 ^ n12955 ;
  assign n13825 = n13817 ^ n12955 ;
  assign n13827 = n13826 ^ n13825 ;
  assign n13828 = n13816 & ~n13827 ;
  assign n13829 = n13828 ^ n13826 ;
  assign n13831 = n13830 ^ n13829 ;
  assign n13832 = n13831 ^ n12955 ;
  assign n13833 = ~n12420 & n13832 ;
  assign n13834 = n13833 ^ n12955 ;
  assign n13850 = n13849 ^ n13834 ;
  assign n13959 = n13850 ^ x337 ;
  assign n13958 = n13952 ^ n13850 ;
  assign n13960 = n13959 ^ n13958 ;
  assign n13961 = n13957 & ~n13960 ;
  assign n13962 = n13961 ^ n13959 ;
  assign n14054 = n13962 ^ x336 ;
  assign n14133 = n14091 ^ n14054 ;
  assign n14264 = n13471 & ~n14133 ;
  assign n14265 = n14264 ^ n13472 ;
  assign n14346 = n14265 ^ n12735 ;
  assign n14347 = x487 & n14346 ;
  assign n14266 = n12735 & n14265 ;
  assign n14344 = n14266 ^ n12737 ;
  assign n14092 = ~n14054 & ~n14091 ;
  assign n13851 = n13850 ^ x336 ;
  assign n13963 = ~n13851 & n13962 ;
  assign n13964 = n13963 ^ x336 ;
  assign n14052 = n13964 ^ x351 ;
  assign n13845 = n12947 ^ n12943 ;
  assign n13840 = n13830 ^ n12955 ;
  assign n13841 = n13829 & n13840 ;
  assign n13842 = n13841 ^ n12955 ;
  assign n13839 = n13415 ^ n13414 ;
  assign n13843 = n13842 ^ n13839 ;
  assign n13844 = ~n12946 & n13843 ;
  assign n13846 = n13845 ^ n13844 ;
  assign n13847 = n13846 ^ n11779 ;
  assign n13835 = n13834 ^ n13824 ;
  assign n13836 = n13834 ^ n11768 ;
  assign n13837 = ~n13835 & n13836 ;
  assign n13838 = n13837 ^ n11768 ;
  assign n13848 = n13847 ^ n13838 ;
  assign n14053 = n14052 ^ n13848 ;
  assign n14136 = n14092 ^ n14053 ;
  assign n14135 = n14133 & n14134 ;
  assign n14137 = n14136 ^ n14135 ;
  assign n14267 = ~n13474 & ~n14137 ;
  assign n14138 = n13476 ^ n13475 ;
  assign n14268 = n14267 ^ n14138 ;
  assign n14345 = n14344 ^ n14268 ;
  assign n14348 = n14347 ^ n14345 ;
  assign n14269 = n14268 ^ n14266 ;
  assign n14270 = n14268 ^ n12737 ;
  assign n14271 = n14269 & ~n14270 ;
  assign n14272 = n14271 ^ n12737 ;
  assign n14349 = n14272 ^ n12732 ;
  assign n14139 = n14138 ^ n14135 ;
  assign n14140 = ~n14137 & n14139 ;
  assign n14141 = n14140 ^ n14136 ;
  assign n14093 = ~n14053 & n14092 ;
  assign n13965 = n13964 ^ n13848 ;
  assign n13966 = n13846 ^ n13838 ;
  assign n13967 = n13417 ^ n13416 ;
  assign n13968 = n13967 ^ n13845 ;
  assign n13969 = n13968 ^ n13842 ;
  assign n13970 = n13969 ^ n13967 ;
  assign n13971 = ~n13843 & n13970 ;
  assign n13972 = n13971 ^ n13968 ;
  assign n13973 = ~n13120 & ~n13972 ;
  assign n13974 = n13973 ^ n12951 ;
  assign n13975 = n13974 ^ n11779 ;
  assign n13976 = n13975 ^ n13974 ;
  assign n13977 = n13976 ^ n13838 ;
  assign n13978 = ~n13966 & n13977 ;
  assign n13979 = n13978 ^ n13975 ;
  assign n13980 = n13979 ^ n12664 ;
  assign n13981 = n13980 ^ x351 ;
  assign n13982 = n13981 ^ n13848 ;
  assign n13983 = n13982 ^ n13980 ;
  assign n13984 = n13965 & ~n13983 ;
  assign n13985 = n13984 ^ n13981 ;
  assign n14051 = n13985 ^ x350 ;
  assign n14131 = n14093 ^ n14051 ;
  assign n14273 = n14141 ^ n14131 ;
  assign n14274 = n13468 & n14273 ;
  assign n14130 = n13480 ^ n13469 ;
  assign n14275 = n14274 ^ n14130 ;
  assign n14350 = n14349 ^ n14275 ;
  assign n14351 = n14350 ^ x486 ;
  assign n14352 = n14351 ^ n14345 ;
  assign n14353 = n14352 ^ n14350 ;
  assign n14354 = n14348 & ~n14353 ;
  assign n14355 = n14354 ^ n14351 ;
  assign n14276 = n14275 ^ n14272 ;
  assign n14277 = n14275 ^ n12732 ;
  assign n14278 = ~n14276 & n14277 ;
  assign n14279 = n14278 ^ n12732 ;
  assign n14356 = n14279 ^ n12727 ;
  assign n14132 = n14131 ^ n14130 ;
  assign n14142 = n14141 ^ n14130 ;
  assign n14143 = ~n14132 & n14142 ;
  assign n14144 = n14143 ^ n14131 ;
  assign n14094 = ~n14051 & ~n14093 ;
  assign n13998 = n13974 ^ n12664 ;
  assign n13999 = n13979 & ~n13998 ;
  assign n14000 = n13999 ^ n12664 ;
  assign n14001 = n14000 ^ n11966 ;
  assign n13993 = n13419 ^ n13418 ;
  assign n13987 = n13127 ^ n12670 ;
  assign n13989 = n13987 ^ n13967 ;
  assign n13986 = n13120 ^ n12951 ;
  assign n13988 = n13987 ^ n13986 ;
  assign n13990 = n13989 ^ n13988 ;
  assign n13991 = n13972 & n13990 ;
  assign n13992 = n13991 ^ n13989 ;
  assign n13994 = n13993 ^ n13992 ;
  assign n13995 = n13994 ^ n13127 ;
  assign n13996 = n12670 & ~n13995 ;
  assign n13997 = n13996 ^ n13994 ;
  assign n14002 = n14001 ^ n13997 ;
  assign n14004 = n14002 ^ x350 ;
  assign n14003 = n14002 ^ n13980 ;
  assign n14005 = n14004 ^ n14003 ;
  assign n14006 = ~n13985 & n14005 ;
  assign n14007 = n14006 ^ n14004 ;
  assign n14050 = n14007 ^ x349 ;
  assign n14128 = n14094 ^ n14050 ;
  assign n14280 = n14144 ^ n14128 ;
  assign n14281 = ~n13465 & n14280 ;
  assign n14126 = n13482 ^ n13465 ;
  assign n14127 = n14126 ^ n13464 ;
  assign n14282 = n14281 ^ n14127 ;
  assign n14357 = n14356 ^ n14282 ;
  assign n14359 = n14357 ^ x485 ;
  assign n14358 = n14357 ^ n14350 ;
  assign n14360 = n14359 ^ n14358 ;
  assign n14361 = ~n14355 & n14360 ;
  assign n14362 = n14361 ^ n14359 ;
  assign n14283 = n14282 ^ n14279 ;
  assign n14284 = n14282 ^ n12727 ;
  assign n14285 = n14283 & ~n14284 ;
  assign n14286 = n14285 ^ n12727 ;
  assign n14363 = n14286 ^ n12724 ;
  assign n14129 = n14128 ^ n14127 ;
  assign n14145 = n14144 ^ n14127 ;
  assign n14146 = n14129 & ~n14145 ;
  assign n14147 = n14146 ^ n14128 ;
  assign n14095 = n14050 & ~n14094 ;
  assign n14014 = n13993 ^ n13987 ;
  assign n14015 = n13992 & n14014 ;
  assign n14013 = n13987 ^ n13302 ;
  assign n14016 = n14015 ^ n14013 ;
  assign n14012 = n13421 ^ n13420 ;
  assign n14017 = n14016 ^ n14012 ;
  assign n14018 = n14017 ^ n13302 ;
  assign n14019 = ~n12791 & n14018 ;
  assign n14020 = n14019 ^ n13302 ;
  assign n14008 = n14000 ^ n13997 ;
  assign n14009 = ~n14001 & ~n14008 ;
  assign n14010 = n14009 ^ n11966 ;
  assign n14011 = n14010 ^ n12784 ;
  assign n14021 = n14020 ^ n14011 ;
  assign n14023 = n14021 ^ x349 ;
  assign n14022 = n14021 ^ n14002 ;
  assign n14024 = n14023 ^ n14022 ;
  assign n14025 = ~n14007 & n14024 ;
  assign n14026 = n14025 ^ n14023 ;
  assign n14049 = n14026 ^ x348 ;
  assign n14125 = n14095 ^ n14049 ;
  assign n14148 = n14147 ^ n14125 ;
  assign n14261 = n13461 & n14148 ;
  assign n14149 = n13485 ^ n13461 ;
  assign n14150 = n14149 ^ n13459 ;
  assign n14262 = n14261 ^ n14150 ;
  assign n14364 = n14363 ^ n14262 ;
  assign n14366 = n14364 ^ x484 ;
  assign n14365 = n14364 ^ n14357 ;
  assign n14367 = n14366 ^ n14365 ;
  assign n14368 = n14362 & ~n14367 ;
  assign n14369 = n14368 ^ n14366 ;
  assign n14151 = n14150 ^ n14125 ;
  assign n14152 = n14148 & n14151 ;
  assign n14153 = n14152 ^ n14147 ;
  assign n14096 = ~n14049 & n14095 ;
  assign n14037 = n13423 ^ n13422 ;
  assign n14032 = n13323 ^ n13302 ;
  assign n14033 = n14032 ^ n13323 ;
  assign n14034 = n14033 ^ n14012 ;
  assign n14035 = n14016 & n14034 ;
  assign n14036 = n14035 ^ n14032 ;
  assign n14038 = n14037 ^ n14036 ;
  assign n14039 = n14038 ^ n13323 ;
  assign n14040 = ~n12820 & ~n14039 ;
  assign n14041 = n14040 ^ n13323 ;
  assign n14027 = n14020 ^ n14010 ;
  assign n14028 = n14020 ^ n12784 ;
  assign n14029 = n14027 & ~n14028 ;
  assign n14030 = n14029 ^ n12784 ;
  assign n14031 = n14030 ^ n12006 ;
  assign n14042 = n14041 ^ n14031 ;
  assign n14044 = n14042 ^ x348 ;
  assign n14043 = n14042 ^ n14021 ;
  assign n14045 = n14044 ^ n14043 ;
  assign n14046 = n14026 & ~n14045 ;
  assign n14047 = n14046 ^ n14044 ;
  assign n14048 = n14047 ^ x347 ;
  assign n14123 = n14096 ^ n14048 ;
  assign n14291 = n14153 ^ n14123 ;
  assign n14292 = ~n13489 & ~n14291 ;
  assign n14121 = n13489 ^ n13377 ;
  assign n14122 = n14121 ^ n13488 ;
  assign n14293 = n14292 ^ n14122 ;
  assign n14263 = n14262 ^ n12724 ;
  assign n14287 = n14286 ^ n14262 ;
  assign n14288 = ~n14263 & ~n14287 ;
  assign n14289 = n14288 ^ n12724 ;
  assign n14290 = n14289 ^ n12719 ;
  assign n14370 = n14293 ^ n14290 ;
  assign n14372 = n14370 ^ x483 ;
  assign n14371 = n14370 ^ n14364 ;
  assign n14373 = n14372 ^ n14371 ;
  assign n14374 = n14369 & ~n14373 ;
  assign n14375 = n14374 ^ n14372 ;
  assign n14124 = n14123 ^ n14122 ;
  assign n14154 = n14153 ^ n14122 ;
  assign n14155 = ~n14124 & ~n14154 ;
  assign n14156 = n14155 ^ n14123 ;
  assign n14108 = n13426 ^ n13424 ;
  assign n14104 = n13344 ^ n13323 ;
  assign n14103 = n14037 ^ n13344 ;
  assign n14105 = n14104 ^ n14103 ;
  assign n14106 = n14036 & ~n14105 ;
  assign n14107 = n14106 ^ n14104 ;
  assign n14109 = n14108 ^ n14107 ;
  assign n14110 = n14109 ^ n13344 ;
  assign n14111 = n12840 & ~n14110 ;
  assign n14112 = n14111 ^ n13344 ;
  assign n14098 = n14041 ^ n14030 ;
  assign n14099 = n14041 ^ n12006 ;
  assign n14100 = n14098 & n14099 ;
  assign n14101 = n14100 ^ n12006 ;
  assign n14102 = n14101 ^ n12833 ;
  assign n14113 = n14112 ^ n14102 ;
  assign n14115 = n14113 ^ x347 ;
  assign n14114 = n14113 ^ n14042 ;
  assign n14116 = n14115 ^ n14114 ;
  assign n14117 = ~n14047 & n14116 ;
  assign n14118 = n14117 ^ n14115 ;
  assign n14119 = n14118 ^ x346 ;
  assign n14097 = n14048 & n14096 ;
  assign n14120 = n14119 ^ n14097 ;
  assign n14157 = n14156 ^ n14120 ;
  assign n14298 = ~n13492 & ~n14157 ;
  assign n14299 = n14298 ^ n13697 ;
  assign n14294 = n14293 ^ n14289 ;
  assign n14295 = ~n14290 & ~n14294 ;
  assign n14296 = n14295 ^ n12719 ;
  assign n14297 = n14296 ^ n12716 ;
  assign n14376 = n14299 ^ n14297 ;
  assign n14378 = n14376 ^ x482 ;
  assign n14377 = n14376 ^ n14370 ;
  assign n14379 = n14378 ^ n14377 ;
  assign n14380 = ~n14375 & n14379 ;
  assign n14381 = n14380 ^ n14378 ;
  assign n14183 = n14097 & ~n14119 ;
  assign n14171 = n13428 ^ n13427 ;
  assign n14167 = n13365 ^ n13344 ;
  assign n14166 = n14108 ^ n13365 ;
  assign n14168 = n14167 ^ n14166 ;
  assign n14169 = n14107 & ~n14168 ;
  assign n14170 = n14169 ^ n14167 ;
  assign n14172 = n14171 ^ n14170 ;
  assign n14173 = n14172 ^ n13365 ;
  assign n14174 = ~n12867 & ~n14173 ;
  assign n14175 = n14174 ^ n13365 ;
  assign n14161 = n14112 ^ n14101 ;
  assign n14162 = n14112 ^ n12833 ;
  assign n14163 = ~n14161 & n14162 ;
  assign n14164 = n14163 ^ n12833 ;
  assign n14165 = n14164 ^ n12176 ;
  assign n14176 = n14175 ^ n14165 ;
  assign n14178 = n14176 ^ x346 ;
  assign n14177 = n14176 ^ n14113 ;
  assign n14179 = n14178 ^ n14177 ;
  assign n14180 = n14118 & ~n14179 ;
  assign n14181 = n14180 ^ n14178 ;
  assign n14182 = n14181 ^ x345 ;
  assign n14184 = n14183 ^ n14182 ;
  assign n14158 = n14156 ^ n13697 ;
  assign n14159 = n14157 & n14158 ;
  assign n14160 = n14159 ^ n13697 ;
  assign n14185 = n14184 ^ n14160 ;
  assign n14304 = ~n13500 & n14185 ;
  assign n14305 = n14304 ^ n13693 ;
  assign n14300 = n14299 ^ n14296 ;
  assign n14301 = ~n14297 & ~n14300 ;
  assign n14302 = n14301 ^ n12716 ;
  assign n14303 = n14302 ^ n12712 ;
  assign n14382 = n14305 ^ n14303 ;
  assign n14384 = n14382 ^ x481 ;
  assign n14383 = n14382 ^ n14376 ;
  assign n14385 = n14384 ^ n14383 ;
  assign n14386 = n14381 & ~n14385 ;
  assign n14387 = n14386 ^ n14384 ;
  assign n14207 = n14183 ^ n14176 ;
  assign n14208 = ~n14181 & ~n14207 ;
  assign n14205 = n14183 ^ n14181 ;
  assign n14206 = ~x345 & n14205 ;
  assign n14209 = n14208 ^ n14206 ;
  assign n14199 = n14171 ^ n13365 ;
  assign n14200 = ~n14170 & ~n14199 ;
  assign n14196 = n13430 ^ n13429 ;
  assign n14197 = n14196 ^ n13455 ;
  assign n14198 = n14197 ^ n14171 ;
  assign n14201 = n14200 ^ n14198 ;
  assign n14202 = n14201 ^ n13455 ;
  assign n14203 = ~n12917 & ~n14202 ;
  assign n14193 = n13455 ^ n12206 ;
  assign n14192 = n12176 ^ x344 ;
  assign n14194 = n14193 ^ n14192 ;
  assign n14189 = n14175 ^ n14164 ;
  assign n14190 = n14175 ^ n12176 ;
  assign n14191 = ~n14189 & ~n14190 ;
  assign n14195 = n14194 ^ n14191 ;
  assign n14204 = n14203 ^ n14195 ;
  assign n14210 = n14209 ^ n14204 ;
  assign n14186 = n14184 ^ n13693 ;
  assign n14187 = ~n14185 & ~n14186 ;
  assign n14188 = n14187 ^ n13693 ;
  assign n14211 = n14210 ^ n14188 ;
  assign n14310 = n13508 & n14211 ;
  assign n14311 = n14310 ^ n13688 ;
  assign n14306 = n14305 ^ n14302 ;
  assign n14307 = ~n14303 & ~n14306 ;
  assign n14308 = n14307 ^ n12712 ;
  assign n14309 = n14308 ^ n12708 ;
  assign n14388 = n14311 ^ n14309 ;
  assign n14390 = n14388 ^ x480 ;
  assign n14389 = n14388 ^ n14382 ;
  assign n14391 = n14390 ^ n14389 ;
  assign n14392 = ~n14387 & n14391 ;
  assign n14393 = n14392 ^ n14390 ;
  assign n14212 = n14210 ^ n13688 ;
  assign n14213 = ~n14211 & n14212 ;
  assign n14214 = n14213 ^ n13688 ;
  assign n14215 = n14214 ^ n13630 ;
  assign n14316 = n13516 & ~n14215 ;
  assign n14317 = n14316 ^ n13683 ;
  assign n14312 = n14311 ^ n14308 ;
  assign n14313 = ~n14309 & n14312 ;
  assign n14314 = n14313 ^ n12708 ;
  assign n14315 = n14314 ^ n12704 ;
  assign n14394 = n14317 ^ n14315 ;
  assign n14396 = n14394 ^ x495 ;
  assign n14395 = n14394 ^ n14388 ;
  assign n14397 = n14396 ^ n14395 ;
  assign n14398 = ~n14393 & n14397 ;
  assign n14399 = n14398 ^ n14396 ;
  assign n14537 = n14399 ^ x494 ;
  assign n14538 = n14346 ^ x487 ;
  assign n14539 = n14347 ^ x486 ;
  assign n14540 = n14539 ^ n14345 ;
  assign n14541 = n14538 & ~n14540 ;
  assign n14542 = n14355 ^ x485 ;
  assign n14543 = n14541 & n14542 ;
  assign n14544 = n14362 ^ x484 ;
  assign n14545 = n14543 & ~n14544 ;
  assign n14546 = n14369 ^ x483 ;
  assign n14547 = n14545 & ~n14546 ;
  assign n14548 = n14375 ^ x482 ;
  assign n14549 = n14547 & n14548 ;
  assign n14550 = n14381 ^ x481 ;
  assign n14551 = n14549 & ~n14550 ;
  assign n14552 = n14387 ^ x480 ;
  assign n14553 = ~n14551 & ~n14552 ;
  assign n14554 = n14393 ^ x495 ;
  assign n14555 = ~n14553 & n14554 ;
  assign n14556 = ~n14537 & ~n14555 ;
  assign n14318 = n14317 ^ n14314 ;
  assign n14319 = ~n14315 & ~n14318 ;
  assign n14320 = n14319 ^ n12704 ;
  assign n14400 = n14320 ^ n12700 ;
  assign n14218 = n13683 ^ n13646 ;
  assign n14216 = n13683 ^ n13630 ;
  assign n14217 = n14215 & ~n14216 ;
  assign n14219 = n14218 ^ n14217 ;
  assign n13649 = n13632 ^ n13630 ;
  assign n14256 = n14219 ^ n13649 ;
  assign n14257 = n14256 ^ n13646 ;
  assign n14258 = ~n13524 & n14257 ;
  assign n14259 = n14258 ^ n13646 ;
  assign n14401 = n14400 ^ n14259 ;
  assign n14403 = n14401 ^ x494 ;
  assign n14402 = n14401 ^ n14394 ;
  assign n14404 = n14403 ^ n14402 ;
  assign n14405 = ~n14399 & n14404 ;
  assign n14406 = n14405 ^ n14403 ;
  assign n14557 = n14406 ^ x493 ;
  assign n14558 = n14556 & n14557 ;
  assign n14260 = n14259 ^ n12700 ;
  assign n14321 = n14320 ^ n14259 ;
  assign n14322 = ~n14260 & n14321 ;
  assign n14323 = n14322 ^ n12700 ;
  assign n14407 = n14323 ^ n12696 ;
  assign n14224 = n13633 ^ n13629 ;
  assign n13650 = n13649 ^ n13646 ;
  assign n14220 = n13650 & n14219 ;
  assign n13648 = n13647 ^ n13646 ;
  assign n14221 = n14220 ^ n13648 ;
  assign n14251 = n14224 ^ n14221 ;
  assign n14252 = n14251 ^ n13647 ;
  assign n14253 = n13532 & ~n14252 ;
  assign n14254 = n14253 ^ n13647 ;
  assign n14408 = n14407 ^ n14254 ;
  assign n14410 = n14408 ^ x493 ;
  assign n14409 = n14408 ^ n14401 ;
  assign n14411 = n14410 ^ n14409 ;
  assign n14412 = n14406 & ~n14411 ;
  assign n14413 = n14412 ^ n14410 ;
  assign n14559 = n14413 ^ x492 ;
  assign n14560 = ~n14558 & ~n14559 ;
  assign n14255 = n14254 ^ n12696 ;
  assign n14324 = n14323 ^ n14254 ;
  assign n14325 = ~n14255 & ~n14324 ;
  assign n14326 = n14325 ^ n12696 ;
  assign n14414 = n14326 ^ n12693 ;
  assign n13644 = n13635 ^ n13634 ;
  assign n14222 = n13647 ^ n13644 ;
  assign n14223 = n14222 ^ n13644 ;
  assign n14225 = n14224 ^ n14223 ;
  assign n14226 = ~n14221 & n14225 ;
  assign n14227 = n14226 ^ n14222 ;
  assign n14248 = ~n13539 & n14227 ;
  assign n14249 = n14248 ^ n13641 ;
  assign n14415 = n14414 ^ n14249 ;
  assign n14417 = n14415 ^ x492 ;
  assign n14416 = n14415 ^ n14408 ;
  assign n14418 = n14417 ^ n14416 ;
  assign n14419 = n14413 & ~n14418 ;
  assign n14420 = n14419 ^ n14417 ;
  assign n14561 = n14420 ^ x491 ;
  assign n14562 = n14560 & ~n14561 ;
  assign n14250 = n14249 ^ n12693 ;
  assign n14327 = n14326 ^ n14249 ;
  assign n14328 = n14250 & n14327 ;
  assign n14329 = n14328 ^ n12693 ;
  assign n14421 = n14329 ^ n12689 ;
  assign n14232 = n13637 ^ n13636 ;
  assign n13645 = n13644 ^ n13641 ;
  assign n14228 = n13645 & ~n14227 ;
  assign n13643 = n13642 ^ n13641 ;
  assign n14229 = n14228 ^ n13643 ;
  assign n14243 = n14232 ^ n14229 ;
  assign n14244 = n14243 ^ n13642 ;
  assign n14245 = ~n13546 & n14244 ;
  assign n14246 = n14245 ^ n13642 ;
  assign n14422 = n14421 ^ n14246 ;
  assign n14424 = n14422 ^ x491 ;
  assign n14423 = n14422 ^ n14415 ;
  assign n14425 = n14424 ^ n14423 ;
  assign n14426 = n14420 & ~n14425 ;
  assign n14427 = n14426 ^ n14424 ;
  assign n14563 = n14427 ^ x490 ;
  assign n14564 = ~n14562 & ~n14563 ;
  assign n14233 = n14232 ^ n13642 ;
  assign n14234 = n14229 & n14233 ;
  assign n13560 = n13559 ^ n13558 ;
  assign n14230 = n13642 ^ n13560 ;
  assign n14235 = n14234 ^ n14230 ;
  assign n13639 = n13638 ^ n13628 ;
  assign n14334 = n14235 ^ n13639 ;
  assign n14335 = n14334 ^ n13558 ;
  assign n14336 = n13559 & n14335 ;
  assign n14337 = n14336 ^ n13558 ;
  assign n14247 = n14246 ^ n12689 ;
  assign n14330 = n14329 ^ n14246 ;
  assign n14331 = n14247 & ~n14330 ;
  assign n14332 = n14331 ^ n12689 ;
  assign n14333 = n14332 ^ n12219 ;
  assign n14428 = n14337 ^ n14333 ;
  assign n14430 = n14428 ^ x490 ;
  assign n14429 = n14428 ^ n14422 ;
  assign n14431 = n14430 ^ n14429 ;
  assign n14432 = ~n14427 & n14431 ;
  assign n14433 = n14432 ^ n14430 ;
  assign n14565 = n14433 ^ x489 ;
  assign n14566 = n14564 & n14565 ;
  assign n14338 = n14337 ^ n14332 ;
  assign n14339 = ~n14333 & ~n14338 ;
  assign n14340 = n14339 ^ n12219 ;
  assign n14341 = n14340 ^ n12384 ;
  assign n14238 = n14056 ^ n14055 ;
  assign n13640 = n13639 ^ n13560 ;
  assign n14236 = n13640 & n14235 ;
  assign n13567 = n13566 ^ n13560 ;
  assign n14237 = n14236 ^ n13567 ;
  assign n14239 = n14238 ^ n14237 ;
  assign n14240 = n14239 ^ n13566 ;
  assign n14241 = n12807 & ~n14240 ;
  assign n14242 = n14241 ^ n13566 ;
  assign n14342 = n14341 ^ n14242 ;
  assign n14435 = n14342 ^ x489 ;
  assign n14434 = n14428 ^ n14342 ;
  assign n14436 = n14435 ^ n14434 ;
  assign n14437 = n14433 & ~n14436 ;
  assign n14438 = n14437 ^ n14435 ;
  assign n14567 = n14438 ^ x488 ;
  assign n14568 = n14566 & n14567 ;
  assign n14343 = n14342 ^ x488 ;
  assign n14439 = ~n14343 & n14438 ;
  assign n14440 = n14439 ^ x488 ;
  assign n14569 = n14440 ^ x503 ;
  assign n14451 = n14340 ^ n14242 ;
  assign n14452 = ~n14341 & n14451 ;
  assign n14453 = n14452 ^ n12384 ;
  assign n14447 = n13659 ^ n13656 ;
  assign n14448 = n14447 ^ n13655 ;
  assign n14444 = n14058 ^ n14057 ;
  assign n14441 = n14238 ^ n13566 ;
  assign n14442 = n14237 & ~n14441 ;
  assign n14443 = n14442 ^ n13566 ;
  assign n14445 = n14444 ^ n14443 ;
  assign n14446 = ~n13659 & n14445 ;
  assign n14449 = n14448 ^ n14446 ;
  assign n14450 = n14449 ^ n12884 ;
  assign n14454 = n14453 ^ n14450 ;
  assign n14570 = n14569 ^ n14454 ;
  assign n14571 = n14568 & ~n14570 ;
  assign n14455 = n14454 ^ n14440 ;
  assign n14456 = n14453 ^ n14449 ;
  assign n14466 = n14453 ^ n12884 ;
  assign n14467 = n14456 & ~n14466 ;
  assign n14459 = n14448 ^ n14444 ;
  assign n14460 = ~n14445 & ~n14459 ;
  assign n14457 = n14060 ^ n14059 ;
  assign n14458 = n14457 ^ n14448 ;
  assign n14461 = n14460 ^ n14458 ;
  assign n14462 = n13652 & n14461 ;
  assign n14463 = n14462 ^ n13664 ;
  assign n14464 = n14463 ^ n12884 ;
  assign n14468 = n14467 ^ n14464 ;
  assign n14469 = n14468 ^ n12881 ;
  assign n14470 = n14469 ^ x503 ;
  assign n14471 = n14470 ^ n14440 ;
  assign n14472 = n14471 ^ n14469 ;
  assign n14473 = ~n14455 & n14472 ;
  assign n14474 = n14473 ^ n14470 ;
  assign n14572 = n14474 ^ x502 ;
  assign n14573 = ~n14571 & n14572 ;
  assign n14483 = n14463 ^ n12881 ;
  assign n14484 = n14468 & ~n14483 ;
  assign n14485 = n14484 ^ n12881 ;
  assign n14486 = n14485 ^ n12286 ;
  assign n14477 = n13664 ^ n13652 ;
  assign n14478 = n14477 ^ n14457 ;
  assign n14479 = ~n14461 & n14478 ;
  assign n14475 = n14062 ^ n14061 ;
  assign n14476 = n14475 ^ n14457 ;
  assign n14480 = n14479 ^ n14476 ;
  assign n14481 = n13757 & n14480 ;
  assign n14482 = n14481 ^ n13763 ;
  assign n14487 = n14486 ^ n14482 ;
  assign n14489 = n14487 ^ x502 ;
  assign n14488 = n14487 ^ n14469 ;
  assign n14490 = n14489 ^ n14488 ;
  assign n14491 = ~n14474 & n14490 ;
  assign n14492 = n14491 ^ n14489 ;
  assign n14536 = n14492 ^ x501 ;
  assign n14604 = n14573 ^ n14536 ;
  assign n14647 = n14134 & ~n14604 ;
  assign n14648 = n14647 ^ n14133 ;
  assign n14652 = n14648 ^ n13471 ;
  assign n14653 = x135 & n14652 ;
  assign n14649 = n13471 & n14648 ;
  assign n14650 = n14649 ^ n13474 ;
  assign n14605 = n14134 ^ n14133 ;
  assign n14606 = n14604 & n14605 ;
  assign n14574 = n14536 & n14573 ;
  assign n14503 = n14485 ^ n14482 ;
  assign n14504 = ~n14486 & ~n14503 ;
  assign n14505 = n14504 ^ n12286 ;
  assign n14506 = n14505 ^ n12281 ;
  assign n14495 = n13763 ^ n13757 ;
  assign n14496 = n14495 ^ n14475 ;
  assign n14497 = ~n14480 & n14496 ;
  assign n14494 = n14475 ^ n13778 ;
  assign n14498 = n14497 ^ n14494 ;
  assign n14493 = n14064 ^ n14063 ;
  assign n14499 = n14498 ^ n14493 ;
  assign n14500 = n14499 ^ n13778 ;
  assign n14501 = n13771 & n14500 ;
  assign n14502 = n14501 ^ n13778 ;
  assign n14507 = n14506 ^ n14502 ;
  assign n14509 = n14507 ^ x501 ;
  assign n14508 = n14507 ^ n14487 ;
  assign n14510 = n14509 ^ n14508 ;
  assign n14511 = ~n14492 & n14510 ;
  assign n14512 = n14511 ^ n14509 ;
  assign n14535 = n14512 ^ x500 ;
  assign n14603 = n14574 ^ n14535 ;
  assign n14607 = n14606 ^ n14603 ;
  assign n14645 = ~n14138 & ~n14607 ;
  assign n14608 = n14139 ^ n14136 ;
  assign n14646 = n14645 ^ n14608 ;
  assign n14651 = n14650 ^ n14646 ;
  assign n14654 = n14653 ^ n14651 ;
  assign n14609 = n14608 ^ n14603 ;
  assign n14610 = ~n14607 & n14609 ;
  assign n14611 = n14610 ^ n14606 ;
  assign n14575 = ~n14535 & n14574 ;
  assign n14524 = n14505 ^ n14502 ;
  assign n14525 = ~n14506 & ~n14524 ;
  assign n14526 = n14525 ^ n12281 ;
  assign n14527 = n14526 ^ n12276 ;
  assign n14519 = n14066 ^ n14065 ;
  assign n14513 = n13791 ^ n13081 ;
  assign n14514 = n14513 ^ n13778 ;
  assign n14515 = n14514 ^ n14513 ;
  assign n14516 = n14515 ^ n14493 ;
  assign n14517 = ~n14498 & ~n14516 ;
  assign n14518 = n14517 ^ n14514 ;
  assign n14520 = n14519 ^ n14518 ;
  assign n14521 = n14520 ^ n13791 ;
  assign n14522 = n13081 & ~n14521 ;
  assign n14523 = n14522 ^ n14520 ;
  assign n14528 = n14527 ^ n14523 ;
  assign n14530 = n14528 ^ x500 ;
  assign n14529 = n14528 ^ n14507 ;
  assign n14531 = n14530 ^ n14529 ;
  assign n14532 = n14512 & ~n14531 ;
  assign n14533 = n14532 ^ n14530 ;
  assign n14534 = n14533 ^ x499 ;
  assign n14600 = n14575 ^ n14534 ;
  assign n14612 = n14611 ^ n14600 ;
  assign n14659 = n14130 & ~n14612 ;
  assign n14601 = n14142 ^ n14131 ;
  assign n14660 = n14659 ^ n14601 ;
  assign n14655 = n14649 ^ n14646 ;
  assign n14656 = ~n14650 & ~n14655 ;
  assign n14657 = n14656 ^ n13474 ;
  assign n14658 = n14657 ^ n13468 ;
  assign n14661 = n14660 ^ n14658 ;
  assign n14662 = n14661 ^ x134 ;
  assign n14663 = n14662 ^ n14651 ;
  assign n14664 = n14663 ^ n14661 ;
  assign n14665 = n14654 & ~n14664 ;
  assign n14666 = n14665 ^ n14662 ;
  assign n14602 = n14601 ^ n14600 ;
  assign n14613 = ~n14602 & n14612 ;
  assign n14614 = n14613 ^ n14601 ;
  assign n14586 = n14526 ^ n14523 ;
  assign n14587 = n14527 & ~n14586 ;
  assign n14588 = n14587 ^ n12276 ;
  assign n14589 = n14588 ^ n12271 ;
  assign n14579 = n14519 ^ n14513 ;
  assign n14580 = ~n14518 & ~n14579 ;
  assign n14578 = n14513 ^ n13804 ;
  assign n14581 = n14580 ^ n14578 ;
  assign n14577 = n14068 ^ n14067 ;
  assign n14582 = n14581 ^ n14577 ;
  assign n14583 = n14582 ^ n13804 ;
  assign n14584 = ~n13089 & n14583 ;
  assign n14585 = n14584 ^ n13804 ;
  assign n14590 = n14589 ^ n14585 ;
  assign n14592 = n14590 ^ x499 ;
  assign n14591 = n14590 ^ n14528 ;
  assign n14593 = n14592 ^ n14591 ;
  assign n14594 = n14533 & ~n14593 ;
  assign n14595 = n14594 ^ n14592 ;
  assign n14596 = n14595 ^ x498 ;
  assign n14576 = ~n14534 & n14575 ;
  assign n14597 = n14596 ^ n14576 ;
  assign n14615 = n14614 ^ n14597 ;
  assign n14672 = ~n14127 & ~n14615 ;
  assign n14598 = n14145 ^ n14128 ;
  assign n14673 = n14672 ^ n14598 ;
  assign n14667 = n14660 ^ n14657 ;
  assign n14668 = n14660 ^ n13468 ;
  assign n14669 = n14667 & n14668 ;
  assign n14670 = n14669 ^ n13468 ;
  assign n14671 = n14670 ^ n13465 ;
  assign n14674 = n14673 ^ n14671 ;
  assign n14676 = n14674 ^ x133 ;
  assign n14675 = n14674 ^ n14661 ;
  assign n14677 = n14676 ^ n14675 ;
  assign n14678 = n14666 & ~n14677 ;
  assign n14679 = n14678 ^ n14676 ;
  assign n14632 = n14588 ^ n14585 ;
  assign n14633 = n14589 & n14632 ;
  assign n14634 = n14633 ^ n12271 ;
  assign n14635 = n14634 ^ n12266 ;
  assign n14627 = n14070 ^ n14069 ;
  assign n14622 = n13818 ^ n13804 ;
  assign n14623 = n14622 ^ n13818 ;
  assign n14624 = n14623 ^ n14577 ;
  assign n14625 = ~n14581 & ~n14624 ;
  assign n14626 = n14625 ^ n14622 ;
  assign n14628 = n14627 ^ n14626 ;
  assign n14629 = n14628 ^ n13818 ;
  assign n14630 = ~n13097 & ~n14629 ;
  assign n14631 = n14630 ^ n13818 ;
  assign n14636 = n14635 ^ n14631 ;
  assign n14638 = n14636 ^ x498 ;
  assign n14637 = n14636 ^ n14590 ;
  assign n14639 = n14638 ^ n14637 ;
  assign n14640 = ~n14595 & n14639 ;
  assign n14641 = n14640 ^ n14638 ;
  assign n14642 = n14641 ^ x497 ;
  assign n14621 = ~n14576 & ~n14596 ;
  assign n14643 = n14642 ^ n14621 ;
  assign n14599 = n14598 ^ n14597 ;
  assign n14616 = n14599 & n14615 ;
  assign n14617 = n14616 ^ n14598 ;
  assign n14685 = n14643 ^ n14617 ;
  assign n14686 = n14150 & n14685 ;
  assign n14618 = n14150 ^ n14147 ;
  assign n14619 = n14618 ^ n14125 ;
  assign n14687 = n14686 ^ n14619 ;
  assign n14680 = n14673 ^ n14670 ;
  assign n14681 = n14673 ^ n13465 ;
  assign n14682 = n14680 & n14681 ;
  assign n14683 = n14682 ^ n13465 ;
  assign n14684 = n14683 ^ n13461 ;
  assign n14688 = n14687 ^ n14684 ;
  assign n14690 = n14688 ^ x132 ;
  assign n14689 = n14688 ^ n14674 ;
  assign n14691 = n14690 ^ n14689 ;
  assign n14692 = ~n14679 & n14691 ;
  assign n14693 = n14692 ^ n14690 ;
  assign n15097 = n14693 ^ x131 ;
  assign n15098 = n14679 ^ x132 ;
  assign n15099 = ~n15097 & n15098 ;
  assign n14727 = n14154 ^ n14123 ;
  assign n14713 = n14634 ^ n14631 ;
  assign n14714 = n14635 & n14713 ;
  assign n14715 = n14714 ^ n12266 ;
  assign n14716 = n14715 ^ n12420 ;
  assign n14708 = n14072 ^ n14071 ;
  assign n14704 = n13831 ^ n13818 ;
  assign n14703 = n14627 ^ n13831 ;
  assign n14705 = n14704 ^ n14703 ;
  assign n14706 = n14626 & ~n14705 ;
  assign n14707 = n14706 ^ n14704 ;
  assign n14709 = n14708 ^ n14707 ;
  assign n14710 = n14709 ^ n13831 ;
  assign n14711 = ~n12955 & ~n14710 ;
  assign n14712 = n14711 ^ n13831 ;
  assign n14717 = n14716 ^ n14712 ;
  assign n14719 = n14717 ^ x497 ;
  assign n14718 = n14717 ^ n14636 ;
  assign n14720 = n14719 ^ n14718 ;
  assign n14721 = ~n14641 & n14720 ;
  assign n14722 = n14721 ^ n14719 ;
  assign n14723 = n14722 ^ x496 ;
  assign n14702 = ~n14621 & n14642 ;
  assign n14724 = n14723 ^ n14702 ;
  assign n14699 = n14643 ^ n14619 ;
  assign n14700 = ~n14685 & ~n14699 ;
  assign n14701 = n14700 ^ n14619 ;
  assign n14725 = n14724 ^ n14701 ;
  assign n14726 = ~n14122 & n14725 ;
  assign n14728 = n14727 ^ n14726 ;
  assign n14694 = n14687 ^ n14683 ;
  assign n14695 = n14687 ^ n13461 ;
  assign n14696 = n14694 & n14695 ;
  assign n14697 = n14696 ^ n13461 ;
  assign n14698 = n14697 ^ n13489 ;
  assign n14729 = n14728 ^ n14698 ;
  assign n14731 = n14729 ^ x131 ;
  assign n14730 = n14729 ^ n14688 ;
  assign n14732 = n14731 ^ n14730 ;
  assign n14733 = n14693 & ~n14732 ;
  assign n14734 = n14733 ^ n14731 ;
  assign n15100 = n14734 ^ x130 ;
  assign n15101 = n15099 & ~n15100 ;
  assign n14763 = n14158 ^ n14120 ;
  assign n14751 = n14708 ^ n13831 ;
  assign n14752 = ~n14707 & n14751 ;
  assign n14753 = n14752 ^ n13831 ;
  assign n14750 = n14074 ^ n14073 ;
  assign n14754 = n14753 ^ n14750 ;
  assign n14755 = ~n13845 & ~n14754 ;
  assign n14756 = n14755 ^ n13843 ;
  assign n14757 = n14756 ^ n12946 ;
  assign n14747 = n14715 ^ n14712 ;
  assign n14748 = n14716 & ~n14747 ;
  assign n14749 = n14748 ^ n12420 ;
  assign n14758 = n14757 ^ n14749 ;
  assign n14743 = n14717 ^ x496 ;
  assign n14744 = n14722 & ~n14743 ;
  assign n14745 = n14744 ^ x496 ;
  assign n14746 = n14745 ^ x511 ;
  assign n14759 = n14758 ^ n14746 ;
  assign n14742 = ~n14702 & n14723 ;
  assign n14760 = n14759 ^ n14742 ;
  assign n14739 = n14727 ^ n14724 ;
  assign n14740 = ~n14725 & n14739 ;
  assign n14741 = n14740 ^ n14727 ;
  assign n14761 = n14760 ^ n14741 ;
  assign n14762 = n13697 & ~n14761 ;
  assign n14764 = n14763 ^ n14762 ;
  assign n14735 = n14728 ^ n14697 ;
  assign n14736 = ~n14698 & ~n14735 ;
  assign n14737 = n14736 ^ n13489 ;
  assign n14738 = n14737 ^ n13492 ;
  assign n14765 = n14764 ^ n14738 ;
  assign n14767 = n14765 ^ x130 ;
  assign n14766 = n14765 ^ n14729 ;
  assign n14768 = n14767 ^ n14766 ;
  assign n14769 = n14734 & ~n14768 ;
  assign n14770 = n14769 ^ n14767 ;
  assign n15102 = n14770 ^ x129 ;
  assign n15103 = ~n15101 & n15102 ;
  assign n14804 = n14160 ^ n13693 ;
  assign n14805 = n14804 ^ n14184 ;
  assign n14779 = n14758 ^ n14745 ;
  assign n14780 = n14756 ^ n14749 ;
  assign n14785 = n14077 ^ n14075 ;
  assign n14781 = n13845 ^ n13843 ;
  assign n14782 = n14781 ^ n14750 ;
  assign n14783 = n14754 & ~n14782 ;
  assign n14784 = n14783 ^ n14753 ;
  assign n14786 = n14785 ^ n14784 ;
  assign n14787 = ~n13986 & n14786 ;
  assign n14788 = n14787 ^ n13972 ;
  assign n14789 = n14788 ^ n12946 ;
  assign n14790 = n14789 ^ n14749 ;
  assign n14791 = n14790 ^ n14788 ;
  assign n14792 = n14780 & n14791 ;
  assign n14793 = n14792 ^ n14789 ;
  assign n14794 = n14793 ^ n13120 ;
  assign n14795 = n14794 ^ x511 ;
  assign n14796 = n14795 ^ n14745 ;
  assign n14797 = n14796 ^ n14794 ;
  assign n14798 = ~n14779 & n14797 ;
  assign n14799 = n14798 ^ n14795 ;
  assign n14800 = n14799 ^ x510 ;
  assign n14778 = ~n14742 & n14759 ;
  assign n14801 = n14800 ^ n14778 ;
  assign n14775 = n14763 ^ n14760 ;
  assign n14776 = n14761 & n14775 ;
  assign n14777 = n14776 ^ n14763 ;
  assign n14802 = n14801 ^ n14777 ;
  assign n14803 = ~n13693 & ~n14802 ;
  assign n14806 = n14805 ^ n14803 ;
  assign n14771 = n14764 ^ n14737 ;
  assign n14772 = n14738 & ~n14771 ;
  assign n14773 = n14772 ^ n13492 ;
  assign n14774 = n14773 ^ n13500 ;
  assign n14807 = n14806 ^ n14774 ;
  assign n14809 = n14807 ^ x129 ;
  assign n14808 = n14807 ^ n14765 ;
  assign n14810 = n14809 ^ n14808 ;
  assign n14811 = n14770 & ~n14810 ;
  assign n14812 = n14811 ^ n14809 ;
  assign n15104 = n14812 ^ x128 ;
  assign n15105 = n15103 & n15104 ;
  assign n14845 = n14188 ^ n13688 ;
  assign n14846 = n14845 ^ n14210 ;
  assign n14825 = n13986 ^ n13972 ;
  assign n14826 = n14825 ^ n14784 ;
  assign n14827 = n14079 ^ n14078 ;
  assign n14828 = n14827 ^ n14785 ;
  assign n14829 = n14828 ^ n14827 ;
  assign n14830 = n14829 ^ n14784 ;
  assign n14831 = ~n14826 & ~n14830 ;
  assign n14832 = n14831 ^ n14828 ;
  assign n14833 = ~n13987 & ~n14832 ;
  assign n14834 = n14833 ^ n13994 ;
  assign n14821 = n14788 ^ n13120 ;
  assign n14822 = n14793 & ~n14821 ;
  assign n14823 = n14822 ^ n13120 ;
  assign n14824 = n14823 ^ n12670 ;
  assign n14835 = n14834 ^ n14824 ;
  assign n14837 = n14835 ^ x510 ;
  assign n14836 = n14835 ^ n14794 ;
  assign n14838 = n14837 ^ n14836 ;
  assign n14839 = ~n14799 & n14838 ;
  assign n14840 = n14839 ^ n14837 ;
  assign n14841 = n14840 ^ x509 ;
  assign n14820 = n14778 & n14800 ;
  assign n14842 = n14841 ^ n14820 ;
  assign n14817 = n14805 ^ n14801 ;
  assign n14818 = n14802 & ~n14817 ;
  assign n14819 = n14818 ^ n14805 ;
  assign n14843 = n14842 ^ n14819 ;
  assign n14844 = ~n13688 & n14843 ;
  assign n14847 = n14846 ^ n14844 ;
  assign n14813 = n14806 ^ n14773 ;
  assign n14814 = n14774 & ~n14813 ;
  assign n14815 = n14814 ^ n13500 ;
  assign n14816 = n14815 ^ n13508 ;
  assign n14848 = n14847 ^ n14816 ;
  assign n14850 = n14848 ^ x128 ;
  assign n14849 = n14848 ^ n14807 ;
  assign n14851 = n14850 ^ n14849 ;
  assign n14852 = n14812 & ~n14851 ;
  assign n14853 = n14852 ^ n14850 ;
  assign n15106 = n14853 ^ x143 ;
  assign n15107 = n15105 & ~n15106 ;
  assign n14887 = n14216 ^ n14214 ;
  assign n14872 = n14082 ^ n14080 ;
  assign n14868 = n14017 ^ n13994 ;
  assign n14867 = n14827 ^ n14017 ;
  assign n14869 = n14868 ^ n14867 ;
  assign n14870 = n14832 & n14869 ;
  assign n14871 = n14870 ^ n14868 ;
  assign n14873 = n14872 ^ n14871 ;
  assign n14874 = n14873 ^ n14017 ;
  assign n14875 = ~n13302 & ~n14874 ;
  assign n14876 = n14875 ^ n14017 ;
  assign n14862 = n14834 ^ n14823 ;
  assign n14863 = n14834 ^ n12670 ;
  assign n14864 = ~n14862 & n14863 ;
  assign n14865 = n14864 ^ n12670 ;
  assign n14866 = n14865 ^ n12791 ;
  assign n14877 = n14876 ^ n14866 ;
  assign n14879 = n14877 ^ x509 ;
  assign n14878 = n14877 ^ n14835 ;
  assign n14880 = n14879 ^ n14878 ;
  assign n14881 = n14840 & ~n14880 ;
  assign n14882 = n14881 ^ n14879 ;
  assign n14883 = n14882 ^ x508 ;
  assign n14861 = n14820 & ~n14841 ;
  assign n14884 = n14883 ^ n14861 ;
  assign n14858 = n14846 ^ n14842 ;
  assign n14859 = ~n14843 & n14858 ;
  assign n14860 = n14859 ^ n14846 ;
  assign n14885 = n14884 ^ n14860 ;
  assign n14886 = ~n13683 & ~n14885 ;
  assign n14888 = n14887 ^ n14886 ;
  assign n14854 = n14847 ^ n14815 ;
  assign n14855 = ~n14816 & ~n14854 ;
  assign n14856 = n14855 ^ n13508 ;
  assign n14857 = n14856 ^ n13516 ;
  assign n14889 = n14888 ^ n14857 ;
  assign n14891 = n14889 ^ x143 ;
  assign n14890 = n14889 ^ n14848 ;
  assign n14892 = n14891 ^ n14890 ;
  assign n14893 = ~n14853 & n14892 ;
  assign n14894 = n14893 ^ n14891 ;
  assign n15108 = n14894 ^ x142 ;
  assign n15109 = n15107 & ~n15108 ;
  assign n14913 = n14084 ^ n14083 ;
  assign n14909 = n14038 ^ n14017 ;
  assign n14908 = n14872 ^ n14038 ;
  assign n14910 = n14909 ^ n14908 ;
  assign n14911 = n14871 & ~n14910 ;
  assign n14912 = n14911 ^ n14909 ;
  assign n14914 = n14913 ^ n14912 ;
  assign n14915 = n14914 ^ n14038 ;
  assign n14916 = ~n13323 & ~n14915 ;
  assign n14917 = n14916 ^ n14038 ;
  assign n14903 = n14876 ^ n14865 ;
  assign n14904 = n14876 ^ n12791 ;
  assign n14905 = ~n14903 & n14904 ;
  assign n14906 = n14905 ^ n12791 ;
  assign n14907 = n14906 ^ n12820 ;
  assign n14918 = n14917 ^ n14907 ;
  assign n14920 = n14918 ^ x508 ;
  assign n14919 = n14918 ^ n14877 ;
  assign n14921 = n14920 ^ n14919 ;
  assign n14922 = n14882 & ~n14921 ;
  assign n14923 = n14922 ^ n14920 ;
  assign n14924 = n14923 ^ x507 ;
  assign n14902 = ~n14861 & n14883 ;
  assign n14925 = n14924 ^ n14902 ;
  assign n14899 = n14887 ^ n14884 ;
  assign n14900 = n14885 & n14899 ;
  assign n14901 = n14900 ^ n14887 ;
  assign n14926 = n14925 ^ n14901 ;
  assign n14927 = ~n13646 & n14926 ;
  assign n14928 = n14927 ^ n14256 ;
  assign n14895 = n14888 ^ n14856 ;
  assign n14896 = n14857 & ~n14895 ;
  assign n14897 = n14896 ^ n13516 ;
  assign n14898 = n14897 ^ n13524 ;
  assign n14929 = n14928 ^ n14898 ;
  assign n14931 = n14929 ^ x142 ;
  assign n14930 = n14929 ^ n14889 ;
  assign n14932 = n14931 ^ n14930 ;
  assign n14933 = ~n14894 & n14932 ;
  assign n14934 = n14933 ^ n14931 ;
  assign n15110 = n14934 ^ x141 ;
  assign n15111 = ~n15109 & n15110 ;
  assign n14953 = n14086 ^ n14085 ;
  assign n14949 = n14109 ^ n14038 ;
  assign n14948 = n14913 ^ n14109 ;
  assign n14950 = n14949 ^ n14948 ;
  assign n14951 = ~n14912 & n14950 ;
  assign n14952 = n14951 ^ n14949 ;
  assign n14954 = n14953 ^ n14952 ;
  assign n14955 = n14954 ^ n14109 ;
  assign n14956 = ~n13344 & n14955 ;
  assign n14957 = n14956 ^ n14109 ;
  assign n14943 = n14917 ^ n14906 ;
  assign n14944 = n14917 ^ n12820 ;
  assign n14945 = n14943 & ~n14944 ;
  assign n14946 = n14945 ^ n12820 ;
  assign n14947 = n14946 ^ n12840 ;
  assign n14958 = n14957 ^ n14947 ;
  assign n14960 = n14958 ^ x507 ;
  assign n14959 = n14958 ^ n14918 ;
  assign n14961 = n14960 ^ n14959 ;
  assign n14962 = ~n14923 & n14961 ;
  assign n14963 = n14962 ^ n14960 ;
  assign n14964 = n14963 ^ x506 ;
  assign n14942 = n14902 & ~n14924 ;
  assign n14965 = n14964 ^ n14942 ;
  assign n14939 = n14925 ^ n14256 ;
  assign n14940 = ~n14926 & ~n14939 ;
  assign n14941 = n14940 ^ n14256 ;
  assign n14966 = n14965 ^ n14941 ;
  assign n14967 = n13647 & ~n14966 ;
  assign n14968 = n14967 ^ n14251 ;
  assign n14935 = n14928 ^ n14897 ;
  assign n14936 = ~n14898 & n14935 ;
  assign n14937 = n14936 ^ n13524 ;
  assign n14938 = n14937 ^ n13532 ;
  assign n14969 = n14968 ^ n14938 ;
  assign n14971 = n14969 ^ x141 ;
  assign n14970 = n14969 ^ n14929 ;
  assign n14972 = n14971 ^ n14970 ;
  assign n14973 = ~n14934 & n14972 ;
  assign n14974 = n14973 ^ n14971 ;
  assign n15112 = n14974 ^ x140 ;
  assign n15113 = ~n15111 & ~n15112 ;
  assign n15003 = n14965 ^ n14251 ;
  assign n15004 = n14966 & ~n15003 ;
  assign n15005 = n15004 ^ n14251 ;
  assign n15001 = ~n14942 & ~n14964 ;
  assign n14989 = n14088 ^ n14087 ;
  assign n14985 = n14172 ^ n14109 ;
  assign n14984 = n14953 ^ n14172 ;
  assign n14986 = n14985 ^ n14984 ;
  assign n14987 = n14952 & n14986 ;
  assign n14988 = n14987 ^ n14985 ;
  assign n14990 = n14989 ^ n14988 ;
  assign n14991 = n14990 ^ n14172 ;
  assign n14992 = ~n13365 & ~n14991 ;
  assign n14993 = n14992 ^ n14172 ;
  assign n14979 = n14957 ^ n14946 ;
  assign n14980 = n14957 ^ n12840 ;
  assign n14981 = n14979 & n14980 ;
  assign n14982 = n14981 ^ n12840 ;
  assign n14983 = n14982 ^ n12867 ;
  assign n14994 = n14993 ^ n14983 ;
  assign n14996 = n14994 ^ x506 ;
  assign n14995 = n14994 ^ n14958 ;
  assign n14997 = n14996 ^ n14995 ;
  assign n14998 = n14963 & ~n14997 ;
  assign n14999 = n14998 ^ n14996 ;
  assign n15000 = n14999 ^ x505 ;
  assign n15002 = n15001 ^ n15000 ;
  assign n15006 = n15005 ^ n15002 ;
  assign n15007 = n13641 & n15006 ;
  assign n15008 = n15007 ^ n14227 ;
  assign n14975 = n14968 ^ n14937 ;
  assign n14976 = ~n14938 & ~n14975 ;
  assign n14977 = n14976 ^ n13532 ;
  assign n14978 = n14977 ^ n13539 ;
  assign n15009 = n15008 ^ n14978 ;
  assign n15011 = n15009 ^ x140 ;
  assign n15010 = n15009 ^ n14969 ;
  assign n15012 = n15011 ^ n15010 ;
  assign n15013 = ~n14974 & n15012 ;
  assign n15014 = n15013 ^ n15011 ;
  assign n15096 = n15014 ^ x139 ;
  assign n15149 = n15113 ^ n15096 ;
  assign n15148 = n14605 ^ n14604 ;
  assign n16142 = n15149 ^ n15148 ;
  assign n15082 = n14540 ^ n14538 ;
  assign n15039 = n14989 ^ n14172 ;
  assign n15040 = ~n14988 & ~n15039 ;
  assign n15036 = n14090 ^ n14089 ;
  assign n15037 = n15036 ^ n14201 ;
  assign n15038 = n15037 ^ n14989 ;
  assign n15041 = n15040 ^ n15038 ;
  assign n15042 = n15041 ^ n14201 ;
  assign n15043 = ~n13455 & ~n15042 ;
  assign n15033 = n14201 ^ n12917 ;
  assign n15032 = n12867 ^ x504 ;
  assign n15034 = n15033 ^ n15032 ;
  assign n15029 = n14993 ^ n14982 ;
  assign n15030 = n14993 ^ n12867 ;
  assign n15031 = ~n15029 & ~n15030 ;
  assign n15035 = n15034 ^ n15031 ;
  assign n15044 = n15043 ^ n15035 ;
  assign n15024 = n15001 ^ n14994 ;
  assign n15027 = n14999 & n15024 ;
  assign n15023 = n14999 ^ n14994 ;
  assign n15025 = n15024 ^ n15023 ;
  assign n15026 = x505 & n15025 ;
  assign n15028 = n15027 ^ n15026 ;
  assign n15045 = n15044 ^ n15028 ;
  assign n15019 = n14227 ^ n13641 ;
  assign n15020 = n15019 ^ n15002 ;
  assign n15021 = ~n15006 & ~n15020 ;
  assign n15022 = n15021 ^ n15005 ;
  assign n15046 = n15045 ^ n15022 ;
  assign n15055 = n15045 ^ n14243 ;
  assign n15056 = n15046 & n15055 ;
  assign n15057 = n15056 ^ n14243 ;
  assign n15058 = n15057 ^ n14538 ;
  assign n15076 = n15057 ^ n14334 ;
  assign n15080 = ~n15058 & ~n15076 ;
  assign n15077 = n14538 ^ n14239 ;
  assign n15081 = n15080 ^ n15077 ;
  assign n15083 = n15082 ^ n15081 ;
  assign n15192 = n14605 & n15149 ;
  assign n15193 = n15192 ^ n14604 ;
  assign n15194 = n15193 ^ n14134 ;
  assign n15776 = x295 & n15194 ;
  assign n15114 = n15096 & n15113 ;
  assign n15047 = n13642 & ~n15046 ;
  assign n15048 = n15047 ^ n14243 ;
  assign n15015 = n15008 ^ n14977 ;
  assign n15016 = ~n14978 & ~n15015 ;
  assign n15017 = n15016 ^ n13539 ;
  assign n15018 = n15017 ^ n13546 ;
  assign n15049 = n15048 ^ n15018 ;
  assign n15051 = n15049 ^ x139 ;
  assign n15050 = n15049 ^ n15009 ;
  assign n15052 = n15051 ^ n15050 ;
  assign n15053 = n15014 & ~n15052 ;
  assign n15054 = n15053 ^ n15051 ;
  assign n15095 = n15054 ^ x138 ;
  assign n15154 = n15114 ^ n15095 ;
  assign n15150 = n15148 & ~n15149 ;
  assign n15155 = n15154 ^ n15150 ;
  assign n15638 = n14608 & n15155 ;
  assign n15151 = n14608 ^ n14606 ;
  assign n15152 = n15151 ^ n14603 ;
  assign n15639 = n15638 ^ n15152 ;
  assign n15636 = n14134 & n15193 ;
  assign n15637 = n15636 ^ n14138 ;
  assign n15775 = n15639 ^ n15637 ;
  assign n15777 = n15776 ^ n15775 ;
  assign n15153 = n15152 ^ n15150 ;
  assign n15156 = ~n15153 & ~n15155 ;
  assign n15157 = n15156 ^ n15152 ;
  assign n15115 = ~n15095 & n15114 ;
  assign n15061 = n15048 ^ n13546 ;
  assign n15062 = n15048 ^ n15017 ;
  assign n15063 = ~n15061 & n15062 ;
  assign n15064 = n15063 ^ n13546 ;
  assign n15065 = n15064 ^ n13559 ;
  assign n15059 = n13560 & ~n15058 ;
  assign n15060 = n15059 ^ n14334 ;
  assign n15066 = n15065 ^ n15060 ;
  assign n15068 = n15066 ^ x138 ;
  assign n15067 = n15066 ^ n15049 ;
  assign n15069 = n15068 ^ n15067 ;
  assign n15070 = ~n15054 & n15069 ;
  assign n15071 = n15070 ^ n15068 ;
  assign n15094 = n15071 ^ x137 ;
  assign n15146 = n15115 ^ n15094 ;
  assign n15644 = n15157 ^ n15146 ;
  assign n15645 = n14601 & n15644 ;
  assign n15144 = n14611 ^ n14601 ;
  assign n15145 = n15144 ^ n14600 ;
  assign n15646 = n15645 ^ n15145 ;
  assign n15640 = n15639 ^ n15636 ;
  assign n15641 = ~n15637 & n15640 ;
  assign n15642 = n15641 ^ n14138 ;
  assign n15643 = n15642 ^ n14130 ;
  assign n15778 = n15646 ^ n15643 ;
  assign n15779 = n15778 ^ x294 ;
  assign n15780 = n15779 ^ n15775 ;
  assign n15781 = n15780 ^ n15778 ;
  assign n15782 = ~n15777 & n15781 ;
  assign n15783 = n15782 ^ n15779 ;
  assign n15147 = n15146 ^ n15145 ;
  assign n15158 = n15157 ^ n15145 ;
  assign n15159 = n15147 & ~n15158 ;
  assign n15160 = n15159 ^ n15146 ;
  assign n15116 = n15094 & n15115 ;
  assign n15084 = n15083 ^ n14239 ;
  assign n15085 = n13566 & n15084 ;
  assign n15086 = n15085 ^ n14239 ;
  assign n15072 = n15064 ^ n15060 ;
  assign n15073 = ~n15065 & n15072 ;
  assign n15074 = n15073 ^ n13559 ;
  assign n15075 = n15074 ^ n12807 ;
  assign n15087 = n15086 ^ n15075 ;
  assign n15089 = n15087 ^ x137 ;
  assign n15088 = n15087 ^ n15066 ;
  assign n15090 = n15089 ^ n15088 ;
  assign n15091 = n15071 & ~n15090 ;
  assign n15092 = n15091 ^ n15089 ;
  assign n15093 = n15092 ^ x136 ;
  assign n15140 = n15116 ^ n15093 ;
  assign n15161 = n15160 ^ n15140 ;
  assign n15651 = ~n14598 & n15161 ;
  assign n15141 = n14614 ^ n14598 ;
  assign n15142 = n15141 ^ n14597 ;
  assign n15652 = n15651 ^ n15142 ;
  assign n15647 = n15646 ^ n15642 ;
  assign n15648 = ~n15643 & ~n15647 ;
  assign n15649 = n15648 ^ n14130 ;
  assign n15650 = n15649 ^ n14127 ;
  assign n15784 = n15652 ^ n15650 ;
  assign n15786 = n15784 ^ x293 ;
  assign n15785 = n15784 ^ n15778 ;
  assign n15787 = n15786 ^ n15785 ;
  assign n15788 = ~n15783 & n15787 ;
  assign n15789 = n15788 ^ n15786 ;
  assign n15143 = n15142 ^ n15140 ;
  assign n15162 = ~n15143 & ~n15161 ;
  assign n15163 = n15162 ^ n15142 ;
  assign n15122 = n15086 ^ n15074 ;
  assign n15129 = n14459 ^ n14443 ;
  assign n15126 = n14542 ^ n14541 ;
  assign n15123 = n15082 ^ n14239 ;
  assign n15124 = ~n15081 & n15123 ;
  assign n15125 = n15124 ^ n15082 ;
  assign n15127 = n15126 ^ n15125 ;
  assign n15128 = ~n14448 & ~n15127 ;
  assign n15130 = n15129 ^ n15128 ;
  assign n15131 = n15130 ^ n12807 ;
  assign n15132 = n15131 ^ n15130 ;
  assign n15133 = n15132 ^ n15074 ;
  assign n15134 = n15122 & n15133 ;
  assign n15135 = n15134 ^ n15131 ;
  assign n15136 = n15135 ^ n13659 ;
  assign n15118 = n15087 ^ x136 ;
  assign n15119 = n15092 & ~n15118 ;
  assign n15120 = n15119 ^ x136 ;
  assign n15121 = n15120 ^ x151 ;
  assign n15137 = n15136 ^ n15121 ;
  assign n15117 = n15093 & n15116 ;
  assign n15138 = n15137 ^ n15117 ;
  assign n15657 = n15163 ^ n15138 ;
  assign n15658 = n14619 & n15657 ;
  assign n14620 = n14619 ^ n14617 ;
  assign n14644 = n14643 ^ n14620 ;
  assign n15659 = n15658 ^ n14644 ;
  assign n15653 = n15652 ^ n15649 ;
  assign n15654 = ~n15650 & ~n15653 ;
  assign n15655 = n15654 ^ n14127 ;
  assign n15656 = n15655 ^ n14150 ;
  assign n15790 = n15659 ^ n15656 ;
  assign n15792 = n15790 ^ x292 ;
  assign n15791 = n15790 ^ n15784 ;
  assign n15793 = n15792 ^ n15791 ;
  assign n15794 = n15789 & ~n15793 ;
  assign n15795 = n15794 ^ n15792 ;
  assign n15171 = n15136 ^ n15120 ;
  assign n15179 = n15130 ^ n13659 ;
  assign n15180 = n15135 & n15179 ;
  assign n15181 = n15180 ^ n13659 ;
  assign n15182 = n15181 ^ n13652 ;
  assign n15174 = n15129 ^ n15126 ;
  assign n15175 = n15127 & ~n15174 ;
  assign n15172 = n14544 ^ n14543 ;
  assign n15173 = n15172 ^ n15129 ;
  assign n15176 = n15175 ^ n15173 ;
  assign n15177 = n14477 & ~n15176 ;
  assign n15178 = n15177 ^ n14461 ;
  assign n15183 = n15182 ^ n15178 ;
  assign n15184 = n15183 ^ x151 ;
  assign n15185 = n15184 ^ n15120 ;
  assign n15186 = n15185 ^ n15183 ;
  assign n15187 = ~n15171 & n15186 ;
  assign n15188 = n15187 ^ n15184 ;
  assign n15189 = n15188 ^ x150 ;
  assign n15170 = n15117 & ~n15137 ;
  assign n15190 = n15189 ^ n15170 ;
  assign n15139 = n15138 ^ n14644 ;
  assign n15164 = n15163 ^ n14644 ;
  assign n15165 = n15139 & ~n15164 ;
  assign n15166 = n15165 ^ n15138 ;
  assign n15664 = n15190 ^ n15166 ;
  assign n15665 = n14727 & n15664 ;
  assign n15167 = n14727 ^ n14701 ;
  assign n15168 = n15167 ^ n14724 ;
  assign n15666 = n15665 ^ n15168 ;
  assign n15660 = n15659 ^ n15655 ;
  assign n15661 = ~n15656 & n15660 ;
  assign n15662 = n15661 ^ n14150 ;
  assign n15663 = n15662 ^ n14122 ;
  assign n15796 = n15666 ^ n15663 ;
  assign n15798 = n15796 ^ x291 ;
  assign n15797 = n15796 ^ n15790 ;
  assign n15799 = n15798 ^ n15797 ;
  assign n15800 = n15795 & ~n15799 ;
  assign n15801 = n15800 ^ n15798 ;
  assign n15169 = n15168 ^ n15166 ;
  assign n15551 = n15190 ^ n15168 ;
  assign n15552 = ~n15169 & n15551 ;
  assign n15553 = n15552 ^ n15190 ;
  assign n15484 = n15170 & ~n15189 ;
  assign n15257 = n15181 ^ n15178 ;
  assign n15197 = n14495 ^ n14480 ;
  assign n15203 = n15197 ^ n15172 ;
  assign n15200 = n14477 ^ n14461 ;
  assign n15201 = n15200 ^ n15172 ;
  assign n15202 = n15176 & n15201 ;
  assign n15204 = n15203 ^ n15202 ;
  assign n15198 = n14546 ^ n14545 ;
  assign n15252 = n15204 ^ n15198 ;
  assign n15253 = n15252 ^ n14480 ;
  assign n15254 = n14495 & ~n15253 ;
  assign n15255 = n15254 ^ n15252 ;
  assign n15258 = n15255 ^ n13652 ;
  assign n15259 = n15258 ^ n15255 ;
  assign n15260 = n15259 ^ n15178 ;
  assign n15261 = ~n15257 & ~n15260 ;
  assign n15262 = n15261 ^ n15258 ;
  assign n15394 = n15262 ^ n13757 ;
  assign n15396 = n15394 ^ x150 ;
  assign n15395 = n15394 ^ n15183 ;
  assign n15397 = n15396 ^ n15395 ;
  assign n15398 = ~n15188 & n15397 ;
  assign n15399 = n15398 ^ n15396 ;
  assign n15483 = n15399 ^ x149 ;
  assign n15547 = n15484 ^ n15483 ;
  assign n15554 = n15553 ^ n15547 ;
  assign n15671 = ~n14763 & ~n15554 ;
  assign n15548 = n14763 ^ n14741 ;
  assign n15549 = n15548 ^ n14760 ;
  assign n15672 = n15671 ^ n15549 ;
  assign n15667 = n15666 ^ n15662 ;
  assign n15668 = ~n15663 & ~n15667 ;
  assign n15669 = n15668 ^ n14122 ;
  assign n15670 = n15669 ^ n13697 ;
  assign n15802 = n15672 ^ n15670 ;
  assign n15804 = n15802 ^ x290 ;
  assign n15803 = n15802 ^ n15796 ;
  assign n15805 = n15804 ^ n15803 ;
  assign n15806 = n15801 & ~n15805 ;
  assign n15807 = n15806 ^ n15804 ;
  assign n15550 = n15549 ^ n15547 ;
  assign n15555 = ~n15550 & n15554 ;
  assign n15556 = n15555 ^ n15549 ;
  assign n15485 = n15483 & ~n15484 ;
  assign n15207 = n14548 ^ n14547 ;
  assign n15199 = n15198 ^ n15197 ;
  assign n15205 = ~n15199 & n15204 ;
  assign n15206 = n15205 ^ n15198 ;
  assign n15208 = n15207 ^ n15206 ;
  assign n15266 = n13778 & ~n15208 ;
  assign n15267 = n15266 ^ n14499 ;
  assign n15256 = n15255 ^ n13757 ;
  assign n15263 = n15256 & ~n15262 ;
  assign n15264 = n15263 ^ n13757 ;
  assign n15265 = n15264 ^ n13771 ;
  assign n15400 = n15267 ^ n15265 ;
  assign n15402 = n15400 ^ x149 ;
  assign n15401 = n15400 ^ n15394 ;
  assign n15403 = n15402 ^ n15401 ;
  assign n15404 = ~n15399 & n15403 ;
  assign n15405 = n15404 ^ n15402 ;
  assign n15482 = n15405 ^ x148 ;
  assign n15543 = n15485 ^ n15482 ;
  assign n15557 = n15556 ^ n15543 ;
  assign n15677 = ~n14805 & n15557 ;
  assign n15544 = n14805 ^ n14777 ;
  assign n15545 = n15544 ^ n14801 ;
  assign n15678 = n15677 ^ n15545 ;
  assign n15673 = n15672 ^ n15669 ;
  assign n15674 = ~n15670 & n15673 ;
  assign n15675 = n15674 ^ n13697 ;
  assign n15676 = n15675 ^ n13693 ;
  assign n15808 = n15678 ^ n15676 ;
  assign n15810 = n15808 ^ x289 ;
  assign n15809 = n15808 ^ n15802 ;
  assign n15811 = n15810 ^ n15809 ;
  assign n15812 = n15807 & ~n15811 ;
  assign n15813 = n15812 ^ n15810 ;
  assign n15546 = n15545 ^ n15543 ;
  assign n15558 = n15546 & ~n15557 ;
  assign n15559 = n15558 ^ n15545 ;
  assign n15486 = n15482 & n15485 ;
  assign n15214 = n14550 ^ n14549 ;
  assign n15209 = n14520 ^ n14499 ;
  assign n15210 = n15209 ^ n14520 ;
  assign n15211 = n15210 ^ n15206 ;
  assign n15212 = n15208 & ~n15211 ;
  assign n15213 = n15212 ^ n15209 ;
  assign n15272 = n15214 ^ n15213 ;
  assign n15273 = n15272 ^ n14520 ;
  assign n15274 = ~n14513 & ~n15273 ;
  assign n15275 = n15274 ^ n14520 ;
  assign n15268 = n15267 ^ n15264 ;
  assign n15269 = n15265 & ~n15268 ;
  assign n15270 = n15269 ^ n13771 ;
  assign n15271 = n15270 ^ n13081 ;
  assign n15406 = n15275 ^ n15271 ;
  assign n15408 = n15406 ^ x148 ;
  assign n15407 = n15406 ^ n15400 ;
  assign n15409 = n15408 ^ n15407 ;
  assign n15410 = ~n15405 & n15409 ;
  assign n15411 = n15410 ^ n15408 ;
  assign n15481 = n15411 ^ x147 ;
  assign n15541 = n15486 ^ n15481 ;
  assign n15683 = n15559 ^ n15541 ;
  assign n15684 = ~n14846 & ~n15683 ;
  assign n15539 = n14846 ^ n14819 ;
  assign n15540 = n15539 ^ n14842 ;
  assign n15685 = n15684 ^ n15540 ;
  assign n15679 = n15678 ^ n15675 ;
  assign n15680 = ~n15676 & ~n15679 ;
  assign n15681 = n15680 ^ n13693 ;
  assign n15682 = n15681 ^ n13688 ;
  assign n15814 = n15685 ^ n15682 ;
  assign n15816 = n15814 ^ x288 ;
  assign n15815 = n15814 ^ n15808 ;
  assign n15817 = n15816 ^ n15815 ;
  assign n15818 = n15813 & ~n15817 ;
  assign n15819 = n15818 ^ n15816 ;
  assign n15542 = n15541 ^ n15540 ;
  assign n15560 = n15559 ^ n15540 ;
  assign n15561 = n15542 & n15560 ;
  assign n15562 = n15561 ^ n15541 ;
  assign n15487 = ~n15481 & ~n15486 ;
  assign n15220 = n14552 ^ n14551 ;
  assign n15216 = n14582 ^ n14520 ;
  assign n15215 = n15214 ^ n14582 ;
  assign n15217 = n15216 ^ n15215 ;
  assign n15218 = ~n15213 & n15217 ;
  assign n15219 = n15218 ^ n15216 ;
  assign n15280 = n15220 ^ n15219 ;
  assign n15281 = n15280 ^ n14582 ;
  assign n15282 = n13804 & n15281 ;
  assign n15283 = n15282 ^ n14582 ;
  assign n15276 = n15275 ^ n15270 ;
  assign n15277 = ~n15271 & n15276 ;
  assign n15278 = n15277 ^ n13081 ;
  assign n15279 = n15278 ^ n13089 ;
  assign n15412 = n15283 ^ n15279 ;
  assign n15414 = n15412 ^ x147 ;
  assign n15413 = n15412 ^ n15406 ;
  assign n15415 = n15414 ^ n15413 ;
  assign n15416 = ~n15411 & n15415 ;
  assign n15417 = n15416 ^ n15414 ;
  assign n15480 = n15417 ^ x146 ;
  assign n15535 = n15487 ^ n15480 ;
  assign n15563 = n15562 ^ n15535 ;
  assign n15690 = n14887 & n15563 ;
  assign n15536 = n14887 ^ n14860 ;
  assign n15537 = n15536 ^ n14884 ;
  assign n15691 = n15690 ^ n15537 ;
  assign n15686 = n15685 ^ n15681 ;
  assign n15687 = n15682 & ~n15686 ;
  assign n15688 = n15687 ^ n13688 ;
  assign n15689 = n15688 ^ n13683 ;
  assign n15820 = n15691 ^ n15689 ;
  assign n15822 = n15820 ^ x303 ;
  assign n15821 = n15820 ^ n15814 ;
  assign n15823 = n15822 ^ n15821 ;
  assign n15824 = n15819 & ~n15823 ;
  assign n15825 = n15824 ^ n15822 ;
  assign n15538 = n15537 ^ n15535 ;
  assign n15564 = n15538 & ~n15563 ;
  assign n15565 = n15564 ^ n15537 ;
  assign n15488 = n15480 & ~n15487 ;
  assign n15226 = n14554 ^ n14553 ;
  assign n15222 = n14628 ^ n14582 ;
  assign n15221 = n15220 ^ n14628 ;
  assign n15223 = n15222 ^ n15221 ;
  assign n15224 = ~n15219 & ~n15223 ;
  assign n15225 = n15224 ^ n15222 ;
  assign n15227 = n15226 ^ n15225 ;
  assign n15288 = n15227 ^ n14628 ;
  assign n15289 = n13818 & ~n15288 ;
  assign n15290 = n15289 ^ n14628 ;
  assign n15284 = n15283 ^ n15278 ;
  assign n15285 = n15279 & n15284 ;
  assign n15286 = n15285 ^ n13089 ;
  assign n15287 = n15286 ^ n13097 ;
  assign n15418 = n15290 ^ n15287 ;
  assign n15420 = n15418 ^ x146 ;
  assign n15419 = n15418 ^ n15412 ;
  assign n15421 = n15420 ^ n15419 ;
  assign n15422 = ~n15417 & n15421 ;
  assign n15423 = n15422 ^ n15420 ;
  assign n15479 = n15423 ^ x145 ;
  assign n15533 = n15488 ^ n15479 ;
  assign n15696 = n15565 ^ n15533 ;
  assign n15697 = ~n14256 & ~n15696 ;
  assign n15531 = n14901 ^ n14256 ;
  assign n15532 = n15531 ^ n14925 ;
  assign n15698 = n15697 ^ n15532 ;
  assign n15692 = n15691 ^ n15688 ;
  assign n15693 = n15689 & ~n15692 ;
  assign n15694 = n15693 ^ n13683 ;
  assign n15695 = n15694 ^ n13646 ;
  assign n15826 = n15698 ^ n15695 ;
  assign n15828 = n15826 ^ x302 ;
  assign n15827 = n15826 ^ n15820 ;
  assign n15829 = n15828 ^ n15827 ;
  assign n15830 = n15825 & ~n15829 ;
  assign n15831 = n15830 ^ n15828 ;
  assign n16069 = n15831 ^ x301 ;
  assign n16051 = n15776 ^ x294 ;
  assign n16052 = n16051 ^ n15775 ;
  assign n16053 = n15783 ^ x293 ;
  assign n16054 = ~n16052 & ~n16053 ;
  assign n16055 = n15789 ^ x292 ;
  assign n16056 = ~n16054 & ~n16055 ;
  assign n16057 = n15795 ^ x291 ;
  assign n16058 = n16056 & ~n16057 ;
  assign n16059 = n15801 ^ x290 ;
  assign n16060 = ~n16058 & n16059 ;
  assign n16061 = n15807 ^ x289 ;
  assign n16062 = n16060 & n16061 ;
  assign n16063 = n15813 ^ x288 ;
  assign n16064 = n16062 & n16063 ;
  assign n16065 = n15819 ^ x303 ;
  assign n16066 = n16064 & n16065 ;
  assign n16067 = n15825 ^ x302 ;
  assign n16068 = ~n16066 & ~n16067 ;
  assign n16372 = n16069 ^ n16068 ;
  assign n16163 = n15553 ^ n15549 ;
  assign n16164 = n16163 ^ n15547 ;
  assign n15195 = n15194 ^ x295 ;
  assign n15191 = n15190 ^ n15169 ;
  assign n15196 = n15195 ^ n15191 ;
  assign n16132 = n15164 ^ n15138 ;
  assign n16159 = n16132 ^ n15191 ;
  assign n15310 = n14825 ^ n14786 ;
  assign n15244 = n14559 ^ n14558 ;
  assign n15231 = n14557 ^ n14556 ;
  assign n15230 = n14782 ^ n14753 ;
  assign n15232 = n15231 ^ n15230 ;
  assign n15233 = n14555 ^ n14537 ;
  assign n15234 = n15233 ^ n14709 ;
  assign n15237 = n14709 ^ n14628 ;
  assign n15235 = n15226 ^ n14628 ;
  assign n15236 = ~n15225 & n15235 ;
  assign n15238 = n15237 ^ n15236 ;
  assign n15239 = ~n15234 & n15238 ;
  assign n15240 = n15239 ^ n15233 ;
  assign n15241 = n15240 ^ n15230 ;
  assign n15242 = n15232 & ~n15241 ;
  assign n15243 = n15242 ^ n15231 ;
  assign n15245 = n15244 ^ n15243 ;
  assign n15943 = n15310 ^ n15245 ;
  assign n15916 = n15098 ^ n15097 ;
  assign n15295 = n15238 ^ n15233 ;
  assign n15912 = n15295 ^ n15098 ;
  assign n15228 = n14666 ^ x133 ;
  assign n15229 = n15228 ^ n15227 ;
  assign n15612 = n15280 ^ n15227 ;
  assign n15507 = n15208 ^ n14499 ;
  assign n15600 = n15507 ^ n15272 ;
  assign n15249 = n15240 ^ n15231 ;
  assign n15250 = ~n14781 & n15249 ;
  assign n15251 = n15250 ^ n15230 ;
  assign n15431 = n15251 ^ n13845 ;
  assign n15291 = n15290 ^ n15286 ;
  assign n15292 = n15287 & ~n15291 ;
  assign n15293 = n15292 ^ n13097 ;
  assign n15294 = n15293 ^ n12955 ;
  assign n15296 = n15295 ^ n14709 ;
  assign n15297 = ~n13831 & n15296 ;
  assign n15298 = n15297 ^ n14709 ;
  assign n15299 = n15298 ^ n15293 ;
  assign n15300 = n15294 & n15299 ;
  assign n15301 = n15300 ^ n12955 ;
  assign n15432 = n15431 ^ n15301 ;
  assign n15392 = n15298 ^ n15294 ;
  assign n15393 = n15392 ^ x144 ;
  assign n15425 = n15392 ^ x145 ;
  assign n15424 = n15418 ^ n15392 ;
  assign n15426 = n15425 ^ n15424 ;
  assign n15427 = n15423 & ~n15426 ;
  assign n15428 = n15427 ^ n15425 ;
  assign n15429 = n15393 & ~n15428 ;
  assign n15430 = n15429 ^ x144 ;
  assign n15433 = n15432 ^ n15430 ;
  assign n15302 = n15301 ^ n15251 ;
  assign n15246 = ~n14825 & n15245 ;
  assign n15247 = n15246 ^ n14786 ;
  assign n15303 = n15247 ^ n13845 ;
  assign n15304 = n15303 ^ n15251 ;
  assign n15305 = n15304 ^ n15247 ;
  assign n15306 = ~n15302 & n15305 ;
  assign n15307 = n15306 ^ n15303 ;
  assign n15434 = n15307 ^ n13986 ;
  assign n15435 = n15434 ^ x159 ;
  assign n15436 = n15435 ^ n15430 ;
  assign n15437 = n15436 ^ n15434 ;
  assign n15438 = n15433 & n15437 ;
  assign n15439 = n15438 ^ n15435 ;
  assign n15248 = n15247 ^ n13986 ;
  assign n15308 = n15248 & ~n15307 ;
  assign n15309 = n15308 ^ n13986 ;
  assign n15440 = n15309 ^ n13987 ;
  assign n15311 = n15310 ^ n15243 ;
  assign n15312 = n14561 ^ n14560 ;
  assign n15313 = n15312 ^ n15244 ;
  assign n15314 = n15313 ^ n15312 ;
  assign n15315 = n15314 ^ n15243 ;
  assign n15316 = n15311 & ~n15315 ;
  assign n15317 = n15316 ^ n15313 ;
  assign n15318 = ~n13994 & n15317 ;
  assign n15319 = n15318 ^ n14832 ;
  assign n15441 = n15440 ^ n15319 ;
  assign n15443 = n15441 ^ x158 ;
  assign n15442 = n15441 ^ n15434 ;
  assign n15444 = n15443 ^ n15442 ;
  assign n15445 = n15439 & ~n15444 ;
  assign n15446 = n15445 ^ n15443 ;
  assign n15320 = n15319 ^ n15309 ;
  assign n15321 = n15319 ^ n13987 ;
  assign n15322 = ~n15320 & n15321 ;
  assign n15323 = n15322 ^ n13987 ;
  assign n15447 = n15323 ^ n13302 ;
  assign n15329 = n14563 ^ n14562 ;
  assign n15325 = n14832 ^ n13994 ;
  assign n15326 = n15325 ^ n15312 ;
  assign n15327 = ~n15317 & ~n15326 ;
  assign n15324 = n15312 ^ n14873 ;
  assign n15328 = n15327 ^ n15324 ;
  assign n15330 = n15329 ^ n15328 ;
  assign n15331 = n15330 ^ n14873 ;
  assign n15332 = ~n14017 & n15331 ;
  assign n15333 = n15332 ^ n14873 ;
  assign n15448 = n15447 ^ n15333 ;
  assign n15450 = n15448 ^ x157 ;
  assign n15449 = n15448 ^ n15441 ;
  assign n15451 = n15450 ^ n15449 ;
  assign n15452 = n15446 & ~n15451 ;
  assign n15453 = n15452 ^ n15450 ;
  assign n15334 = n15333 ^ n15323 ;
  assign n15335 = n15333 ^ n13302 ;
  assign n15336 = n15334 & ~n15335 ;
  assign n15337 = n15336 ^ n13302 ;
  assign n15454 = n15337 ^ n13323 ;
  assign n15343 = n14565 ^ n14564 ;
  assign n15339 = n14914 ^ n14873 ;
  assign n15338 = n15329 ^ n14914 ;
  assign n15340 = n15339 ^ n15338 ;
  assign n15341 = ~n15328 & ~n15340 ;
  assign n15342 = n15341 ^ n15339 ;
  assign n15344 = n15343 ^ n15342 ;
  assign n15345 = n15344 ^ n14914 ;
  assign n15346 = n14038 & ~n15345 ;
  assign n15347 = n15346 ^ n14914 ;
  assign n15455 = n15454 ^ n15347 ;
  assign n15457 = n15455 ^ x156 ;
  assign n15456 = n15455 ^ n15448 ;
  assign n15458 = n15457 ^ n15456 ;
  assign n15459 = ~n15453 & n15458 ;
  assign n15460 = n15459 ^ n15457 ;
  assign n15348 = n15347 ^ n15337 ;
  assign n15349 = n15347 ^ n13323 ;
  assign n15350 = ~n15348 & n15349 ;
  assign n15351 = n15350 ^ n13323 ;
  assign n15461 = n15351 ^ n13344 ;
  assign n15357 = n14567 ^ n14566 ;
  assign n15353 = n14954 ^ n14914 ;
  assign n15352 = n15343 ^ n14954 ;
  assign n15354 = n15353 ^ n15352 ;
  assign n15355 = ~n15342 & n15354 ;
  assign n15356 = n15355 ^ n15353 ;
  assign n15358 = n15357 ^ n15356 ;
  assign n15359 = n15358 ^ n14954 ;
  assign n15360 = n14109 & n15359 ;
  assign n15361 = n15360 ^ n14954 ;
  assign n15462 = n15461 ^ n15361 ;
  assign n15464 = n15462 ^ x155 ;
  assign n15463 = n15462 ^ n15455 ;
  assign n15465 = n15464 ^ n15463 ;
  assign n15466 = n15460 & ~n15465 ;
  assign n15467 = n15466 ^ n15464 ;
  assign n15362 = n15361 ^ n15351 ;
  assign n15363 = n15361 ^ n13344 ;
  assign n15364 = n15362 & ~n15363 ;
  assign n15365 = n15364 ^ n13344 ;
  assign n15468 = n15365 ^ n13365 ;
  assign n15371 = n14570 ^ n14568 ;
  assign n15367 = n14990 ^ n14954 ;
  assign n15366 = n15357 ^ n14990 ;
  assign n15368 = n15367 ^ n15366 ;
  assign n15369 = ~n15356 & ~n15368 ;
  assign n15370 = n15369 ^ n15367 ;
  assign n15372 = n15371 ^ n15370 ;
  assign n15373 = n15372 ^ n14990 ;
  assign n15374 = n14172 & n15373 ;
  assign n15375 = n15374 ^ n14990 ;
  assign n15469 = n15468 ^ n15375 ;
  assign n15471 = n15469 ^ x154 ;
  assign n15470 = n15469 ^ n15462 ;
  assign n15472 = n15471 ^ n15470 ;
  assign n15473 = ~n15467 & n15472 ;
  assign n15474 = n15473 ^ n15471 ;
  assign n15475 = n15439 ^ x158 ;
  assign n15476 = n15430 ^ x159 ;
  assign n15477 = n15476 ^ n15432 ;
  assign n15478 = n15428 ^ x144 ;
  assign n15489 = n15479 & ~n15488 ;
  assign n15490 = ~n15478 & n15489 ;
  assign n15491 = n15477 & n15490 ;
  assign n15492 = n15475 & n15491 ;
  assign n15493 = n15446 ^ x157 ;
  assign n15494 = n15492 & n15493 ;
  assign n15495 = n15453 ^ x156 ;
  assign n15496 = ~n15494 & n15495 ;
  assign n15497 = n15460 ^ x155 ;
  assign n15498 = n15496 & ~n15497 ;
  assign n15499 = n15467 ^ x154 ;
  assign n15500 = ~n15498 & ~n15499 ;
  assign n15503 = n15500 ^ n15469 ;
  assign n15504 = n15474 & ~n15503 ;
  assign n15501 = n15500 ^ n15474 ;
  assign n15502 = x153 & ~n15501 ;
  assign n15505 = n15504 ^ n15502 ;
  assign n15386 = n15371 ^ n14990 ;
  assign n15387 = n15370 & ~n15386 ;
  assign n15383 = n14572 ^ n14571 ;
  assign n15384 = n15383 ^ n15041 ;
  assign n15385 = n15384 ^ n15371 ;
  assign n15388 = n15387 ^ n15385 ;
  assign n15389 = n15388 ^ n15041 ;
  assign n15390 = n14201 & ~n15389 ;
  assign n15380 = n15041 ^ n13455 ;
  assign n15379 = n13365 ^ x152 ;
  assign n15381 = n15380 ^ n15379 ;
  assign n15376 = n15375 ^ n15365 ;
  assign n15377 = n15375 ^ n13365 ;
  assign n15378 = ~n15376 & n15377 ;
  assign n15382 = n15381 ^ n15378 ;
  assign n15391 = n15390 ^ n15382 ;
  assign n15506 = n15505 ^ n15391 ;
  assign n15508 = n15507 ^ n15506 ;
  assign n15509 = n15474 ^ x153 ;
  assign n15510 = n15509 ^ n15500 ;
  assign n15511 = n15510 ^ n15252 ;
  assign n15513 = n15499 ^ n15498 ;
  assign n15512 = n15200 ^ n15176 ;
  assign n15514 = n15513 ^ n15512 ;
  assign n15586 = n15129 ^ n15127 ;
  assign n15581 = n15495 ^ n15494 ;
  assign n15517 = n15493 ^ n15492 ;
  assign n15515 = n14538 ^ n14334 ;
  assign n15516 = n15515 ^ n15057 ;
  assign n15518 = n15517 ^ n15516 ;
  assign n15520 = n15022 ^ n14243 ;
  assign n15521 = n15520 ^ n15045 ;
  assign n15519 = n15491 ^ n15475 ;
  assign n15522 = n15521 ^ n15519 ;
  assign n15525 = n15490 ^ n15477 ;
  assign n15523 = n15019 ^ n15005 ;
  assign n15524 = n15523 ^ n15002 ;
  assign n15526 = n15525 ^ n15524 ;
  assign n15528 = n14941 ^ n14251 ;
  assign n15529 = n15528 ^ n14965 ;
  assign n15527 = n15489 ^ n15478 ;
  assign n15530 = n15529 ^ n15527 ;
  assign n15534 = n15533 ^ n15532 ;
  assign n15566 = n15565 ^ n15532 ;
  assign n15567 = ~n15534 & ~n15566 ;
  assign n15568 = n15567 ^ n15533 ;
  assign n15569 = n15568 ^ n15527 ;
  assign n15570 = n15530 & ~n15569 ;
  assign n15571 = n15570 ^ n15529 ;
  assign n15572 = n15571 ^ n15524 ;
  assign n15573 = n15526 & n15572 ;
  assign n15574 = n15573 ^ n15525 ;
  assign n15575 = n15574 ^ n15519 ;
  assign n15576 = n15522 & ~n15575 ;
  assign n15577 = n15576 ^ n15521 ;
  assign n15578 = n15577 ^ n15516 ;
  assign n15579 = n15518 & ~n15578 ;
  assign n15580 = n15579 ^ n15517 ;
  assign n15582 = n15581 ^ n15580 ;
  assign n15583 = n15581 ^ n15083 ;
  assign n15584 = ~n15582 & n15583 ;
  assign n15585 = n15584 ^ n15083 ;
  assign n15587 = n15586 ^ n15585 ;
  assign n15588 = n15497 ^ n15496 ;
  assign n15589 = n15588 ^ n15585 ;
  assign n15590 = ~n15587 & ~n15589 ;
  assign n15591 = n15590 ^ n15586 ;
  assign n15592 = n15591 ^ n15512 ;
  assign n15593 = n15514 & n15592 ;
  assign n15594 = n15593 ^ n15513 ;
  assign n15595 = n15594 ^ n15510 ;
  assign n15596 = ~n15511 & ~n15595 ;
  assign n15597 = n15596 ^ n15252 ;
  assign n15598 = n15597 ^ n15506 ;
  assign n15599 = n15508 & n15598 ;
  assign n15601 = n15600 ^ n15599 ;
  assign n15604 = n15280 ^ n15272 ;
  assign n15602 = n14652 ^ x135 ;
  assign n15603 = n15602 ^ n15280 ;
  assign n15605 = n15604 ^ n15603 ;
  assign n15606 = ~n15601 & n15605 ;
  assign n15607 = n15606 ^ n15604 ;
  assign n15608 = n14653 ^ x134 ;
  assign n15609 = n15608 ^ n14651 ;
  assign n15610 = n15609 ^ n15280 ;
  assign n15611 = n15607 & ~n15610 ;
  assign n15613 = n15612 ^ n15611 ;
  assign n15614 = ~n15229 & ~n15613 ;
  assign n15615 = n15614 ^ n15228 ;
  assign n15913 = n15615 ^ n15295 ;
  assign n15914 = ~n15912 & n15913 ;
  assign n15915 = n15914 ^ n15098 ;
  assign n15917 = n15916 ^ n15915 ;
  assign n15919 = n15240 ^ n15232 ;
  assign n15925 = n15919 ^ n15916 ;
  assign n15926 = ~n15917 & n15925 ;
  assign n15927 = n15926 ^ n15919 ;
  assign n15944 = n15943 ^ n15927 ;
  assign n15945 = n15325 ^ n15317 ;
  assign n15928 = n15100 ^ n15099 ;
  assign n15946 = n15945 ^ n15928 ;
  assign n15947 = n15946 ^ n15945 ;
  assign n15948 = n15947 ^ n15927 ;
  assign n15949 = ~n15944 & n15948 ;
  assign n15950 = n15949 ^ n15946 ;
  assign n15951 = n15102 ^ n15101 ;
  assign n15973 = n15951 ^ n15945 ;
  assign n15974 = n15950 & ~n15973 ;
  assign n15972 = n15945 ^ n15330 ;
  assign n15975 = n15974 ^ n15972 ;
  assign n15991 = n15344 ^ n15330 ;
  assign n15992 = n15991 ^ n15344 ;
  assign n15971 = n15104 ^ n15103 ;
  assign n15993 = n15992 ^ n15971 ;
  assign n15994 = ~n15975 & ~n15993 ;
  assign n15995 = n15994 ^ n15991 ;
  assign n16013 = n15358 ^ n15344 ;
  assign n15996 = n15106 ^ n15105 ;
  assign n16012 = n15996 ^ n15358 ;
  assign n16014 = n16013 ^ n16012 ;
  assign n16015 = n15995 & n16014 ;
  assign n16016 = n16015 ^ n16013 ;
  assign n16034 = n15372 ^ n15358 ;
  assign n16017 = n15108 ^ n15107 ;
  assign n16033 = n16017 ^ n15372 ;
  assign n16035 = n16034 ^ n16033 ;
  assign n16036 = n16016 & n16035 ;
  assign n16037 = n16036 ^ n16034 ;
  assign n16038 = n15110 ^ n15109 ;
  assign n16125 = n16038 ^ n15372 ;
  assign n16126 = n16037 & n16125 ;
  assign n16122 = n15388 ^ n15111 ;
  assign n16123 = n16122 ^ n15112 ;
  assign n16124 = n16123 ^ n16038 ;
  assign n16127 = n16126 ^ n16124 ;
  assign n16128 = n16127 ^ n15388 ;
  assign n16129 = ~n15041 & n16128 ;
  assign n16119 = n15388 ^ n14201 ;
  assign n16118 = n14172 ^ x312 ;
  assign n16120 = n16119 ^ n16118 ;
  assign n16039 = n16038 ^ n16037 ;
  assign n16040 = n16039 ^ n15372 ;
  assign n16041 = ~n14990 & ~n16040 ;
  assign n16042 = n16041 ^ n15372 ;
  assign n16018 = n16017 ^ n16016 ;
  assign n16019 = n16018 ^ n15358 ;
  assign n16020 = n14954 & n16019 ;
  assign n16021 = n16020 ^ n15358 ;
  assign n15997 = n15996 ^ n15995 ;
  assign n15998 = n15997 ^ n15344 ;
  assign n15999 = ~n14914 & n15998 ;
  assign n16000 = n15999 ^ n15344 ;
  assign n15976 = n15975 ^ n15971 ;
  assign n15977 = n15976 ^ n15330 ;
  assign n15978 = n14873 & n15977 ;
  assign n15979 = n15978 ^ n15330 ;
  assign n15918 = ~n15230 & n15917 ;
  assign n15920 = n15919 ^ n15918 ;
  assign n15619 = n15609 ^ n15607 ;
  assign n15620 = n15619 ^ n15280 ;
  assign n15621 = n14582 & ~n15620 ;
  assign n15622 = n15621 ^ n15280 ;
  assign n15623 = n15622 ^ n13804 ;
  assign n15628 = n15197 & n15595 ;
  assign n15629 = n15628 ^ n15252 ;
  assign n15630 = n15629 ^ n14495 ;
  assign n15631 = ~n15129 & ~n15589 ;
  assign n15632 = n15631 ^ n15127 ;
  assign n15633 = n15632 ^ n14448 ;
  assign n15699 = n15698 ^ n15694 ;
  assign n15700 = n15695 & ~n15699 ;
  assign n15701 = n15700 ^ n13646 ;
  assign n15702 = n15701 ^ n13647 ;
  assign n15703 = ~n14251 & n15569 ;
  assign n15704 = n15703 ^ n15529 ;
  assign n15705 = n15704 ^ n15701 ;
  assign n15706 = ~n15702 & n15705 ;
  assign n15707 = n15706 ^ n13647 ;
  assign n15708 = n15707 ^ n13641 ;
  assign n15709 = n15571 ^ n15525 ;
  assign n15710 = n15019 & ~n15709 ;
  assign n15711 = n15710 ^ n15524 ;
  assign n15712 = n15711 ^ n15707 ;
  assign n15713 = n15708 & n15712 ;
  assign n15714 = n15713 ^ n13641 ;
  assign n15715 = n15714 ^ n13642 ;
  assign n15716 = n14243 & n15575 ;
  assign n15717 = n15716 ^ n15521 ;
  assign n15718 = n15717 ^ n15714 ;
  assign n15719 = n15715 & n15718 ;
  assign n15720 = n15719 ^ n13642 ;
  assign n15721 = n15720 ^ n13560 ;
  assign n15722 = n15577 ^ n15517 ;
  assign n15723 = n14334 & n15722 ;
  assign n15724 = n15723 ^ n15516 ;
  assign n15725 = n15724 ^ n15720 ;
  assign n15726 = n15721 & n15725 ;
  assign n15727 = n15726 ^ n13560 ;
  assign n15634 = ~n14239 & n15582 ;
  assign n15635 = n15634 ^ n15083 ;
  assign n15728 = n15727 ^ n15635 ;
  assign n15729 = n15632 ^ n13566 ;
  assign n15730 = n15729 ^ n15632 ;
  assign n15731 = n15730 ^ n15635 ;
  assign n15732 = n15728 & ~n15731 ;
  assign n15733 = n15732 ^ n15729 ;
  assign n15734 = n15633 & n15733 ;
  assign n15735 = n15734 ^ n14448 ;
  assign n15736 = n15735 ^ n14477 ;
  assign n15737 = n15591 ^ n15513 ;
  assign n15738 = ~n15200 & n15737 ;
  assign n15739 = n15738 ^ n15176 ;
  assign n15740 = n15739 ^ n15735 ;
  assign n15741 = ~n15736 & n15740 ;
  assign n15742 = n15741 ^ n14477 ;
  assign n15743 = n15742 ^ n15629 ;
  assign n15744 = ~n15630 & ~n15743 ;
  assign n15745 = n15744 ^ n14495 ;
  assign n15746 = n15745 ^ n13778 ;
  assign n15747 = n14499 & n15598 ;
  assign n15748 = n15747 ^ n15208 ;
  assign n15749 = n15748 ^ n15745 ;
  assign n15750 = ~n15746 & ~n15749 ;
  assign n15751 = n15750 ^ n13778 ;
  assign n15624 = n15602 ^ n15601 ;
  assign n15625 = n15624 ^ n15272 ;
  assign n15626 = ~n14520 & ~n15625 ;
  assign n15627 = n15626 ^ n15272 ;
  assign n15752 = n15751 ^ n15627 ;
  assign n15753 = n15622 ^ n14513 ;
  assign n15754 = n15753 ^ n15622 ;
  assign n15755 = n15754 ^ n15627 ;
  assign n15756 = ~n15752 & ~n15755 ;
  assign n15757 = n15756 ^ n15753 ;
  assign n15758 = n15623 & n15757 ;
  assign n15759 = n15758 ^ n13804 ;
  assign n15760 = n15759 ^ n13818 ;
  assign n15761 = n15613 ^ n15228 ;
  assign n15762 = n15761 ^ n15227 ;
  assign n15763 = ~n14628 & ~n15762 ;
  assign n15764 = n15763 ^ n15227 ;
  assign n15765 = n15764 ^ n15759 ;
  assign n15766 = n15760 & ~n15765 ;
  assign n15767 = n15766 ^ n13818 ;
  assign n15768 = n15767 ^ n13831 ;
  assign n15616 = n15615 ^ n15098 ;
  assign n15617 = n14709 & n15616 ;
  assign n15618 = n15617 ^ n15295 ;
  assign n15909 = n15767 ^ n15618 ;
  assign n15910 = ~n15768 & ~n15909 ;
  assign n15911 = n15910 ^ n13831 ;
  assign n15924 = n15920 ^ n15911 ;
  assign n15929 = n15928 ^ n15927 ;
  assign n15930 = n15310 & ~n15929 ;
  assign n15931 = n15930 ^ n15245 ;
  assign n15932 = n15931 ^ n14781 ;
  assign n15933 = n15932 ^ n15911 ;
  assign n15934 = n15933 ^ n15931 ;
  assign n15935 = ~n15924 & n15934 ;
  assign n15936 = n15935 ^ n15932 ;
  assign n15952 = n15951 ^ n15950 ;
  assign n15953 = n15952 ^ n15317 ;
  assign n15954 = ~n15325 & ~n15953 ;
  assign n15955 = n15954 ^ n15952 ;
  assign n15956 = n15955 ^ n14825 ;
  assign n15957 = n15956 ^ n15931 ;
  assign n15958 = n15957 ^ n15955 ;
  assign n15959 = ~n15936 & n15958 ;
  assign n15960 = n15959 ^ n15956 ;
  assign n15967 = n15955 ^ n13994 ;
  assign n15968 = n15960 & ~n15967 ;
  assign n15969 = n15968 ^ n13994 ;
  assign n15986 = n15979 ^ n15969 ;
  assign n15987 = n15979 ^ n14017 ;
  assign n15988 = n15986 & ~n15987 ;
  assign n15989 = n15988 ^ n14017 ;
  assign n16007 = n16000 ^ n15989 ;
  assign n16008 = n16000 ^ n14038 ;
  assign n16009 = n16007 & n16008 ;
  assign n16010 = n16009 ^ n14038 ;
  assign n16028 = n16021 ^ n16010 ;
  assign n16029 = n16021 ^ n14109 ;
  assign n16030 = ~n16028 & n16029 ;
  assign n16031 = n16030 ^ n14109 ;
  assign n16115 = n16042 ^ n16031 ;
  assign n16116 = n16042 ^ n14172 ;
  assign n16117 = n16115 & ~n16116 ;
  assign n16121 = n16120 ^ n16117 ;
  assign n16130 = n16129 ^ n16121 ;
  assign n15921 = n15920 ^ n14781 ;
  assign n15922 = n15921 ^ n15911 ;
  assign n15769 = n15768 ^ n15618 ;
  assign n15770 = n15769 ^ x304 ;
  assign n15772 = n15727 ^ n13566 ;
  assign n15773 = n15772 ^ n15635 ;
  assign n15774 = n15773 ^ x296 ;
  assign n15832 = n15704 ^ n15702 ;
  assign n15834 = n15832 ^ x301 ;
  assign n15833 = n15832 ^ n15826 ;
  assign n15835 = n15834 ^ n15833 ;
  assign n15836 = n15831 & ~n15835 ;
  assign n15837 = n15836 ^ n15834 ;
  assign n15838 = n15711 ^ n15708 ;
  assign n15840 = n15838 ^ x300 ;
  assign n15839 = n15838 ^ n15832 ;
  assign n15841 = n15840 ^ n15839 ;
  assign n15842 = n15837 & ~n15841 ;
  assign n15843 = n15842 ^ n15840 ;
  assign n15844 = n15717 ^ n15715 ;
  assign n15846 = n15844 ^ x299 ;
  assign n15845 = n15844 ^ n15838 ;
  assign n15847 = n15846 ^ n15845 ;
  assign n15848 = n15843 & ~n15847 ;
  assign n15849 = n15848 ^ n15846 ;
  assign n15850 = n15724 ^ n15721 ;
  assign n15852 = n15850 ^ x298 ;
  assign n15851 = n15850 ^ n15844 ;
  assign n15853 = n15852 ^ n15851 ;
  assign n15854 = n15849 & ~n15853 ;
  assign n15855 = n15854 ^ n15852 ;
  assign n15857 = n15773 ^ x297 ;
  assign n15856 = n15850 ^ n15773 ;
  assign n15858 = n15857 ^ n15856 ;
  assign n15859 = n15855 & ~n15858 ;
  assign n15860 = n15859 ^ n15857 ;
  assign n15861 = ~n15774 & n15860 ;
  assign n15862 = n15861 ^ x296 ;
  assign n15771 = n15733 ^ n14448 ;
  assign n15863 = n15862 ^ n15771 ;
  assign n15864 = n15739 ^ n15736 ;
  assign n15865 = n15864 ^ x311 ;
  assign n15866 = n15865 ^ n15771 ;
  assign n15867 = n15866 ^ n15864 ;
  assign n15868 = ~n15863 & n15867 ;
  assign n15869 = n15868 ^ n15865 ;
  assign n15870 = n15742 ^ n14495 ;
  assign n15871 = n15870 ^ n15629 ;
  assign n15873 = n15871 ^ x310 ;
  assign n15872 = n15871 ^ n15864 ;
  assign n15874 = n15873 ^ n15872 ;
  assign n15875 = n15869 & ~n15874 ;
  assign n15876 = n15875 ^ n15873 ;
  assign n15877 = n15748 ^ n15746 ;
  assign n15879 = n15877 ^ x309 ;
  assign n15878 = n15877 ^ n15871 ;
  assign n15880 = n15879 ^ n15878 ;
  assign n15881 = n15876 & ~n15880 ;
  assign n15882 = n15881 ^ n15879 ;
  assign n15883 = n15751 ^ n14513 ;
  assign n15884 = n15883 ^ n15627 ;
  assign n15886 = n15884 ^ x308 ;
  assign n15885 = n15884 ^ n15877 ;
  assign n15887 = n15886 ^ n15885 ;
  assign n15888 = ~n15882 & n15887 ;
  assign n15889 = n15888 ^ n15886 ;
  assign n15890 = n15757 ^ n13804 ;
  assign n15892 = n15890 ^ x307 ;
  assign n15891 = n15890 ^ n15884 ;
  assign n15893 = n15892 ^ n15891 ;
  assign n15894 = n15889 & ~n15893 ;
  assign n15895 = n15894 ^ n15892 ;
  assign n15896 = n15764 ^ n15760 ;
  assign n15898 = n15896 ^ x306 ;
  assign n15897 = n15896 ^ n15890 ;
  assign n15899 = n15898 ^ n15897 ;
  assign n15900 = n15895 & ~n15899 ;
  assign n15901 = n15900 ^ n15898 ;
  assign n15903 = n15769 ^ x305 ;
  assign n15902 = n15896 ^ n15769 ;
  assign n15904 = n15903 ^ n15902 ;
  assign n15905 = ~n15901 & n15904 ;
  assign n15906 = n15905 ^ n15903 ;
  assign n15907 = ~n15770 & n15906 ;
  assign n15908 = n15907 ^ x304 ;
  assign n15923 = n15922 ^ n15908 ;
  assign n15937 = n15936 ^ n14825 ;
  assign n15938 = n15937 ^ x319 ;
  assign n15939 = n15938 ^ n15908 ;
  assign n15940 = n15939 ^ n15937 ;
  assign n15941 = n15923 & n15940 ;
  assign n15942 = n15941 ^ n15938 ;
  assign n15961 = n15960 ^ n13994 ;
  assign n15963 = n15961 ^ x318 ;
  assign n15962 = n15961 ^ n15937 ;
  assign n15964 = n15963 ^ n15962 ;
  assign n15965 = n15942 & ~n15964 ;
  assign n15966 = n15965 ^ n15963 ;
  assign n15970 = n15969 ^ n14017 ;
  assign n15980 = n15979 ^ n15970 ;
  assign n15982 = n15980 ^ x317 ;
  assign n15981 = n15980 ^ n15961 ;
  assign n15983 = n15982 ^ n15981 ;
  assign n15984 = ~n15966 & n15983 ;
  assign n15985 = n15984 ^ n15982 ;
  assign n15990 = n15989 ^ n14038 ;
  assign n16001 = n16000 ^ n15990 ;
  assign n16003 = n16001 ^ x316 ;
  assign n16002 = n16001 ^ n15980 ;
  assign n16004 = n16003 ^ n16002 ;
  assign n16005 = ~n15985 & n16004 ;
  assign n16006 = n16005 ^ n16003 ;
  assign n16011 = n16010 ^ n14109 ;
  assign n16022 = n16021 ^ n16011 ;
  assign n16024 = n16022 ^ x315 ;
  assign n16023 = n16022 ^ n16001 ;
  assign n16025 = n16024 ^ n16023 ;
  assign n16026 = n16006 & ~n16025 ;
  assign n16027 = n16026 ^ n16024 ;
  assign n16032 = n16031 ^ n14172 ;
  assign n16043 = n16042 ^ n16032 ;
  assign n16045 = n16043 ^ x314 ;
  assign n16044 = n16043 ^ n16022 ;
  assign n16046 = n16045 ^ n16044 ;
  assign n16047 = ~n16027 & n16046 ;
  assign n16048 = n16047 ^ n16045 ;
  assign n16050 = n16027 ^ x314 ;
  assign n16070 = ~n16068 & n16069 ;
  assign n16071 = n15837 ^ x300 ;
  assign n16072 = n16070 & n16071 ;
  assign n16073 = n15843 ^ x299 ;
  assign n16074 = ~n16072 & ~n16073 ;
  assign n16075 = n15849 ^ x298 ;
  assign n16076 = n16074 & ~n16075 ;
  assign n16077 = n15855 ^ x297 ;
  assign n16078 = ~n16076 & n16077 ;
  assign n16079 = n15860 ^ x296 ;
  assign n16080 = n16078 & n16079 ;
  assign n16081 = n15862 ^ x311 ;
  assign n16082 = n16081 ^ n15771 ;
  assign n16083 = n16080 & ~n16082 ;
  assign n16084 = n15869 ^ x310 ;
  assign n16085 = ~n16083 & ~n16084 ;
  assign n16086 = n15876 ^ x309 ;
  assign n16087 = n16085 & ~n16086 ;
  assign n16088 = n15882 ^ x308 ;
  assign n16089 = n16087 & n16088 ;
  assign n16090 = n15889 ^ x307 ;
  assign n16091 = n16089 & ~n16090 ;
  assign n16092 = n15895 ^ x306 ;
  assign n16093 = ~n16091 & n16092 ;
  assign n16094 = n15901 ^ x305 ;
  assign n16095 = n16093 & ~n16094 ;
  assign n16096 = n15906 ^ x304 ;
  assign n16097 = n16095 & n16096 ;
  assign n16098 = n15908 ^ x319 ;
  assign n16099 = n16098 ^ n15922 ;
  assign n16100 = n16097 & n16099 ;
  assign n16101 = n15942 ^ x318 ;
  assign n16102 = ~n16100 & ~n16101 ;
  assign n16103 = n15966 ^ x317 ;
  assign n16104 = n16102 & n16103 ;
  assign n16105 = n15985 ^ x316 ;
  assign n16106 = n16104 & n16105 ;
  assign n16107 = n16006 ^ x315 ;
  assign n16108 = n16106 & ~n16107 ;
  assign n16109 = ~n16050 & ~n16108 ;
  assign n16110 = n16109 ^ n16043 ;
  assign n16113 = n16048 & ~n16110 ;
  assign n16049 = n16048 ^ n16043 ;
  assign n16111 = n16110 ^ n16049 ;
  assign n16112 = ~x313 & n16111 ;
  assign n16114 = n16113 ^ n16112 ;
  assign n16131 = n16130 ^ n16114 ;
  assign n16133 = n16132 ^ n16131 ;
  assign n16136 = n15160 ^ n15142 ;
  assign n16137 = n16136 ^ n15140 ;
  assign n16134 = n16048 ^ x313 ;
  assign n16135 = n16134 ^ n16109 ;
  assign n16138 = n16137 ^ n16135 ;
  assign n16140 = n16108 ^ n16050 ;
  assign n16139 = n15158 ^ n15146 ;
  assign n16141 = n16140 ^ n16139 ;
  assign n16145 = n15154 ^ n15153 ;
  assign n16143 = n16105 ^ n16104 ;
  assign n16144 = ~n16142 & n16143 ;
  assign n16146 = n16145 ^ n16144 ;
  assign n16147 = n16107 ^ n16106 ;
  assign n16148 = n16147 ^ n16144 ;
  assign n16149 = ~n16146 & n16148 ;
  assign n16150 = n16149 ^ n16145 ;
  assign n16151 = n16150 ^ n16139 ;
  assign n16152 = n16141 & ~n16151 ;
  assign n16153 = n16152 ^ n16140 ;
  assign n16154 = n16153 ^ n16135 ;
  assign n16155 = n16138 & n16154 ;
  assign n16156 = n16155 ^ n16137 ;
  assign n16157 = n16156 ^ n16131 ;
  assign n16158 = ~n16133 & n16157 ;
  assign n16160 = n16159 ^ n16158 ;
  assign n16161 = n15196 & ~n16160 ;
  assign n16162 = n16161 ^ n15195 ;
  assign n16165 = n16164 ^ n16162 ;
  assign n16166 = n15556 ^ n15545 ;
  assign n16167 = n16166 ^ n15543 ;
  assign n16168 = n16167 ^ n16052 ;
  assign n16169 = n16168 ^ n16167 ;
  assign n16170 = n16169 ^ n16162 ;
  assign n16171 = n16165 & ~n16170 ;
  assign n16172 = n16171 ^ n16168 ;
  assign n16174 = n15560 ^ n15541 ;
  assign n16176 = n16174 ^ n16167 ;
  assign n16173 = n16053 ^ n16052 ;
  assign n16175 = n16174 ^ n16173 ;
  assign n16177 = n16176 ^ n16175 ;
  assign n16178 = ~n16172 & ~n16177 ;
  assign n16179 = n16178 ^ n16176 ;
  assign n16181 = n15562 ^ n15537 ;
  assign n16182 = n16181 ^ n15535 ;
  assign n16184 = n16182 ^ n16174 ;
  assign n16180 = n16055 ^ n16054 ;
  assign n16183 = n16182 ^ n16180 ;
  assign n16185 = n16184 ^ n16183 ;
  assign n16186 = n16179 & n16185 ;
  assign n16187 = n16186 ^ n16184 ;
  assign n16189 = n15566 ^ n15533 ;
  assign n16191 = n16189 ^ n16182 ;
  assign n16188 = n16057 ^ n16056 ;
  assign n16190 = n16189 ^ n16188 ;
  assign n16192 = n16191 ^ n16190 ;
  assign n16193 = ~n16187 & n16192 ;
  assign n16194 = n16193 ^ n16191 ;
  assign n16335 = n15568 ^ n15529 ;
  assign n16336 = n16335 ^ n15527 ;
  assign n16338 = n16336 ^ n16189 ;
  assign n16195 = n16059 ^ n16058 ;
  assign n16337 = n16336 ^ n16195 ;
  assign n16339 = n16338 ^ n16337 ;
  assign n16340 = ~n16194 & n16339 ;
  assign n16341 = n16340 ^ n16338 ;
  assign n16343 = n15572 ^ n15525 ;
  assign n16345 = n16343 ^ n16336 ;
  assign n16342 = n16061 ^ n16060 ;
  assign n16344 = n16343 ^ n16342 ;
  assign n16346 = n16345 ^ n16344 ;
  assign n16347 = n16341 & ~n16346 ;
  assign n16348 = n16347 ^ n16345 ;
  assign n16350 = n15574 ^ n15521 ;
  assign n16351 = n16350 ^ n15519 ;
  assign n16353 = n16351 ^ n16343 ;
  assign n16349 = n16063 ^ n16062 ;
  assign n16352 = n16351 ^ n16349 ;
  assign n16354 = n16353 ^ n16352 ;
  assign n16355 = n16348 & ~n16354 ;
  assign n16356 = n16355 ^ n16353 ;
  assign n16358 = n15578 ^ n15517 ;
  assign n16360 = n16358 ^ n16351 ;
  assign n16357 = n16065 ^ n16064 ;
  assign n16359 = n16358 ^ n16357 ;
  assign n16361 = n16360 ^ n16359 ;
  assign n16362 = ~n16356 & n16361 ;
  assign n16363 = n16362 ^ n16360 ;
  assign n16365 = n15580 ^ n15083 ;
  assign n16366 = n16365 ^ n15581 ;
  assign n16368 = n16366 ^ n16358 ;
  assign n16364 = n16067 ^ n16066 ;
  assign n16367 = n16366 ^ n16364 ;
  assign n16369 = n16368 ^ n16367 ;
  assign n16370 = n16363 & ~n16369 ;
  assign n16371 = n16370 ^ n16368 ;
  assign n16396 = n16372 ^ n16371 ;
  assign n16495 = n16396 ^ n16366 ;
  assign n16496 = ~n15083 & ~n16495 ;
  assign n16497 = n16496 ^ n16366 ;
  assign n16395 = n16364 ^ n16363 ;
  assign n16456 = n16395 ^ n16358 ;
  assign n16457 = ~n15516 & ~n16456 ;
  assign n16458 = n16457 ^ n16358 ;
  assign n16459 = n16458 ^ n14334 ;
  assign n16398 = n16357 ^ n16356 ;
  assign n16460 = n16398 ^ n16351 ;
  assign n16461 = ~n15521 & ~n16460 ;
  assign n16462 = n16461 ^ n16351 ;
  assign n16463 = n16462 ^ n14243 ;
  assign n16400 = n16349 ^ n16348 ;
  assign n16464 = n16400 ^ n16343 ;
  assign n16465 = ~n15524 & ~n16464 ;
  assign n16466 = n16465 ^ n16343 ;
  assign n16467 = n16466 ^ n15019 ;
  assign n16402 = n16342 ^ n16341 ;
  assign n16468 = n16402 ^ n16336 ;
  assign n16469 = n15529 & ~n16468 ;
  assign n16470 = n16469 ^ n16336 ;
  assign n16471 = n16470 ^ n14251 ;
  assign n16196 = n16195 ^ n16194 ;
  assign n16472 = n16196 ^ n16189 ;
  assign n16473 = ~n15532 & ~n16472 ;
  assign n16474 = n16473 ^ n16189 ;
  assign n16475 = n16474 ^ n14256 ;
  assign n16307 = n16188 ^ n16187 ;
  assign n16308 = n16307 ^ n16182 ;
  assign n16309 = ~n15537 & ~n16308 ;
  assign n16310 = n16309 ^ n16182 ;
  assign n16476 = n16310 ^ n14887 ;
  assign n16278 = n16173 ^ n16172 ;
  assign n16279 = n16278 ^ n16167 ;
  assign n16280 = n15545 & n16279 ;
  assign n16281 = n16280 ^ n16167 ;
  assign n16292 = n16281 ^ n14805 ;
  assign n16264 = n16162 ^ n16052 ;
  assign n16265 = n15549 & ~n16264 ;
  assign n16266 = n16265 ^ n16164 ;
  assign n16201 = n15148 & ~n16143 ;
  assign n16202 = n16201 ^ n15149 ;
  assign n16203 = n14605 & ~n16202 ;
  assign n16204 = n16203 ^ n14608 ;
  assign n16199 = ~n15152 & ~n16148 ;
  assign n16200 = n16199 ^ n16145 ;
  assign n16212 = n16203 ^ n16200 ;
  assign n16213 = n16204 & n16212 ;
  assign n16214 = n16213 ^ n14608 ;
  assign n16215 = n16214 ^ n14601 ;
  assign n16209 = n16150 ^ n16140 ;
  assign n16210 = ~n15145 & n16209 ;
  assign n16211 = n16210 ^ n16139 ;
  assign n16224 = n16214 ^ n16211 ;
  assign n16225 = n16215 & n16224 ;
  assign n16226 = n16225 ^ n14601 ;
  assign n16227 = n16226 ^ n14598 ;
  assign n16222 = n15142 & ~n16154 ;
  assign n16223 = n16222 ^ n16137 ;
  assign n16236 = n16226 ^ n16223 ;
  assign n16237 = ~n16227 & ~n16236 ;
  assign n16238 = n16237 ^ n14598 ;
  assign n16239 = n16238 ^ n14619 ;
  assign n16234 = n14644 & ~n16157 ;
  assign n16235 = n16234 ^ n16132 ;
  assign n16250 = n16238 ^ n16235 ;
  assign n16251 = ~n16239 & n16250 ;
  assign n16252 = n16251 ^ n14619 ;
  assign n16253 = n16252 ^ n14727 ;
  assign n16246 = n16160 ^ n15195 ;
  assign n16247 = n16246 ^ n15191 ;
  assign n16248 = n15168 & n16247 ;
  assign n16249 = n16248 ^ n15191 ;
  assign n16260 = n16252 ^ n16249 ;
  assign n16261 = n16253 & ~n16260 ;
  assign n16262 = n16261 ^ n14727 ;
  assign n16273 = n16266 ^ n16262 ;
  assign n16274 = n16266 ^ n14763 ;
  assign n16275 = n16273 & n16274 ;
  assign n16276 = n16275 ^ n14763 ;
  assign n16293 = n16281 ^ n16276 ;
  assign n16294 = ~n16292 & n16293 ;
  assign n16295 = n16294 ^ n14805 ;
  assign n16296 = n16295 ^ n14846 ;
  assign n16288 = n16180 ^ n16179 ;
  assign n16289 = n16288 ^ n16174 ;
  assign n16290 = ~n15540 & n16289 ;
  assign n16291 = n16290 ^ n16174 ;
  assign n16303 = n16295 ^ n16291 ;
  assign n16304 = n16296 & n16303 ;
  assign n16305 = n16304 ^ n14846 ;
  assign n16477 = n16310 ^ n16305 ;
  assign n16478 = ~n16476 & ~n16477 ;
  assign n16479 = n16478 ^ n14887 ;
  assign n16480 = n16479 ^ n16474 ;
  assign n16481 = ~n16475 & ~n16480 ;
  assign n16482 = n16481 ^ n14256 ;
  assign n16483 = n16482 ^ n16470 ;
  assign n16484 = ~n16471 & n16483 ;
  assign n16485 = n16484 ^ n14251 ;
  assign n16486 = n16485 ^ n16466 ;
  assign n16487 = n16467 & n16486 ;
  assign n16488 = n16487 ^ n15019 ;
  assign n16489 = n16488 ^ n16462 ;
  assign n16490 = ~n16463 & n16489 ;
  assign n16491 = n16490 ^ n14243 ;
  assign n16492 = n16491 ^ n16458 ;
  assign n16493 = ~n16459 & n16492 ;
  assign n16494 = n16493 ^ n14334 ;
  assign n16498 = n16497 ^ n16494 ;
  assign n16375 = n16071 ^ n16070 ;
  assign n16376 = n16375 ^ n16366 ;
  assign n16373 = n16372 ^ n16366 ;
  assign n16374 = n16371 & ~n16373 ;
  assign n16377 = n16376 ^ n16374 ;
  assign n16499 = n15586 & n16377 ;
  assign n16378 = n15588 ^ n15587 ;
  assign n16500 = n16499 ^ n16378 ;
  assign n16501 = n16500 ^ n14239 ;
  assign n16502 = n16501 ^ n16494 ;
  assign n16503 = n16502 ^ n16500 ;
  assign n16504 = n16498 & ~n16503 ;
  assign n16505 = n16504 ^ n16501 ;
  assign n16587 = n16505 ^ n15129 ;
  assign n16542 = n16494 ^ n14239 ;
  assign n16543 = n16542 ^ n16497 ;
  assign n16544 = n16543 ^ x456 ;
  assign n16206 = n16202 ^ n14605 ;
  assign n16207 = x455 & ~n16206 ;
  assign n16205 = n16204 ^ n16200 ;
  assign n16208 = n16207 ^ n16205 ;
  assign n16216 = n16215 ^ n16211 ;
  assign n16217 = n16216 ^ x454 ;
  assign n16218 = n16217 ^ n16205 ;
  assign n16219 = n16218 ^ n16216 ;
  assign n16220 = n16208 & ~n16219 ;
  assign n16221 = n16220 ^ n16217 ;
  assign n16228 = n16227 ^ n16223 ;
  assign n16230 = n16228 ^ x453 ;
  assign n16229 = n16228 ^ n16216 ;
  assign n16231 = n16230 ^ n16229 ;
  assign n16232 = n16221 & ~n16231 ;
  assign n16233 = n16232 ^ n16230 ;
  assign n16240 = n16239 ^ n16235 ;
  assign n16242 = n16240 ^ x452 ;
  assign n16241 = n16240 ^ n16228 ;
  assign n16243 = n16242 ^ n16241 ;
  assign n16244 = n16233 & ~n16243 ;
  assign n16245 = n16244 ^ n16242 ;
  assign n16254 = n16253 ^ n16249 ;
  assign n16256 = n16254 ^ x451 ;
  assign n16255 = n16254 ^ n16240 ;
  assign n16257 = n16256 ^ n16255 ;
  assign n16258 = n16245 & ~n16257 ;
  assign n16259 = n16258 ^ n16256 ;
  assign n16263 = n16262 ^ n14763 ;
  assign n16267 = n16266 ^ n16263 ;
  assign n16269 = n16267 ^ x450 ;
  assign n16268 = n16267 ^ n16254 ;
  assign n16270 = n16269 ^ n16268 ;
  assign n16271 = ~n16259 & n16270 ;
  assign n16272 = n16271 ^ n16269 ;
  assign n16277 = n16276 ^ n14805 ;
  assign n16282 = n16281 ^ n16277 ;
  assign n16284 = n16282 ^ x449 ;
  assign n16283 = n16282 ^ n16267 ;
  assign n16285 = n16284 ^ n16283 ;
  assign n16286 = ~n16272 & n16285 ;
  assign n16287 = n16286 ^ n16284 ;
  assign n16297 = n16296 ^ n16291 ;
  assign n16299 = n16297 ^ x448 ;
  assign n16298 = n16297 ^ n16282 ;
  assign n16300 = n16299 ^ n16298 ;
  assign n16301 = ~n16287 & n16300 ;
  assign n16302 = n16301 ^ n16299 ;
  assign n16306 = n16305 ^ n14887 ;
  assign n16311 = n16310 ^ n16306 ;
  assign n16313 = n16311 ^ x463 ;
  assign n16312 = n16311 ^ n16297 ;
  assign n16314 = n16313 ^ n16312 ;
  assign n16315 = ~n16302 & n16314 ;
  assign n16316 = n16315 ^ n16313 ;
  assign n16545 = n16479 ^ n14256 ;
  assign n16546 = n16545 ^ n16474 ;
  assign n16548 = n16546 ^ x462 ;
  assign n16547 = n16546 ^ n16311 ;
  assign n16549 = n16548 ^ n16547 ;
  assign n16550 = ~n16316 & n16549 ;
  assign n16551 = n16550 ^ n16548 ;
  assign n16552 = n16482 ^ n14251 ;
  assign n16553 = n16552 ^ n16470 ;
  assign n16555 = n16553 ^ x461 ;
  assign n16554 = n16553 ^ n16546 ;
  assign n16556 = n16555 ^ n16554 ;
  assign n16557 = n16551 & ~n16556 ;
  assign n16558 = n16557 ^ n16555 ;
  assign n16559 = n16485 ^ n15019 ;
  assign n16560 = n16559 ^ n16466 ;
  assign n16562 = n16560 ^ x460 ;
  assign n16561 = n16560 ^ n16553 ;
  assign n16563 = n16562 ^ n16561 ;
  assign n16564 = ~n16558 & n16563 ;
  assign n16565 = n16564 ^ n16562 ;
  assign n16566 = n16488 ^ n14243 ;
  assign n16567 = n16566 ^ n16462 ;
  assign n16569 = n16567 ^ x459 ;
  assign n16568 = n16567 ^ n16560 ;
  assign n16570 = n16569 ^ n16568 ;
  assign n16571 = n16565 & ~n16570 ;
  assign n16572 = n16571 ^ n16569 ;
  assign n16573 = n16491 ^ n14334 ;
  assign n16574 = n16573 ^ n16458 ;
  assign n16576 = n16574 ^ x458 ;
  assign n16575 = n16574 ^ n16567 ;
  assign n16577 = n16576 ^ n16575 ;
  assign n16578 = n16572 & ~n16577 ;
  assign n16579 = n16578 ^ n16576 ;
  assign n16581 = n16543 ^ x457 ;
  assign n16580 = n16574 ^ n16543 ;
  assign n16582 = n16581 ^ n16580 ;
  assign n16583 = n16579 & ~n16582 ;
  assign n16584 = n16583 ^ n16581 ;
  assign n16585 = n16544 & ~n16584 ;
  assign n16586 = n16585 ^ x456 ;
  assign n16588 = n16587 ^ n16586 ;
  assign n16381 = n16073 ^ n16072 ;
  assign n16382 = n16381 ^ n16375 ;
  assign n16379 = n16378 ^ n16375 ;
  assign n16380 = n16377 & ~n16379 ;
  assign n16383 = n16382 ^ n16380 ;
  assign n16453 = ~n15512 & ~n16383 ;
  assign n16384 = n15592 ^ n15513 ;
  assign n16454 = n16453 ^ n16384 ;
  assign n16507 = n16454 ^ n15129 ;
  assign n16506 = n16500 ^ n16454 ;
  assign n16508 = n16507 ^ n16506 ;
  assign n16509 = n16505 & ~n16508 ;
  assign n16510 = n16509 ^ n16507 ;
  assign n16589 = n16510 ^ n15200 ;
  assign n16590 = n16589 ^ x471 ;
  assign n16591 = n16590 ^ n16586 ;
  assign n16592 = n16591 ^ n16589 ;
  assign n16593 = ~n16588 & n16592 ;
  assign n16594 = n16593 ^ n16590 ;
  assign n16455 = n16454 ^ n15200 ;
  assign n16511 = ~n16455 & n16510 ;
  assign n16512 = n16511 ^ n15200 ;
  assign n16595 = n16512 ^ n15197 ;
  assign n16197 = n15594 ^ n15252 ;
  assign n16198 = n16197 ^ n15510 ;
  assign n16389 = n16384 ^ n16198 ;
  assign n16387 = n16384 ^ n16381 ;
  assign n16388 = n16383 & n16387 ;
  assign n16390 = n16389 ^ n16388 ;
  assign n16386 = n16075 ^ n16074 ;
  assign n16391 = n16390 ^ n16386 ;
  assign n16449 = n16391 ^ n16198 ;
  assign n16450 = n15252 & ~n16449 ;
  assign n16451 = n16450 ^ n16198 ;
  assign n16596 = n16595 ^ n16451 ;
  assign n16598 = n16596 ^ x470 ;
  assign n16597 = n16596 ^ n16589 ;
  assign n16599 = n16598 ^ n16597 ;
  assign n16600 = ~n16594 & n16599 ;
  assign n16601 = n16600 ^ n16598 ;
  assign n16452 = n16451 ^ n15197 ;
  assign n16513 = n16512 ^ n16451 ;
  assign n16514 = n16452 & n16513 ;
  assign n16515 = n16514 ^ n15197 ;
  assign n16602 = n16515 ^ n14499 ;
  assign n16406 = n15597 ^ n15507 ;
  assign n16407 = n16406 ^ n15506 ;
  assign n16411 = n16407 ^ n16198 ;
  assign n16412 = n16411 ^ n16407 ;
  assign n16413 = n16412 ^ n16386 ;
  assign n16414 = n16390 & ~n16413 ;
  assign n16415 = n16414 ^ n16411 ;
  assign n16409 = n16077 ^ n16076 ;
  assign n16444 = n16415 ^ n16409 ;
  assign n16445 = n16444 ^ n16407 ;
  assign n16446 = ~n15507 & n16445 ;
  assign n16447 = n16446 ^ n16407 ;
  assign n16603 = n16602 ^ n16447 ;
  assign n16605 = n16603 ^ x469 ;
  assign n16604 = n16603 ^ n16596 ;
  assign n16606 = n16605 ^ n16604 ;
  assign n16607 = n16601 & ~n16606 ;
  assign n16608 = n16607 ^ n16605 ;
  assign n16448 = n16447 ^ n14499 ;
  assign n16516 = n16515 ^ n16447 ;
  assign n16517 = n16448 & ~n16516 ;
  assign n16518 = n16517 ^ n14499 ;
  assign n16609 = n16518 ^ n14520 ;
  assign n16418 = n16079 ^ n16078 ;
  assign n16410 = n16409 ^ n16407 ;
  assign n16416 = n16410 & n16415 ;
  assign n16408 = n16407 ^ n15624 ;
  assign n16417 = n16416 ^ n16408 ;
  assign n16439 = n16418 ^ n16417 ;
  assign n16440 = n16439 ^ n15624 ;
  assign n16441 = n15272 & ~n16440 ;
  assign n16442 = n16441 ^ n15624 ;
  assign n16610 = n16609 ^ n16442 ;
  assign n16612 = n16610 ^ x468 ;
  assign n16611 = n16610 ^ n16603 ;
  assign n16613 = n16612 ^ n16611 ;
  assign n16614 = ~n16608 & n16613 ;
  assign n16615 = n16614 ^ n16612 ;
  assign n16443 = n16442 ^ n14520 ;
  assign n16519 = n16518 ^ n16442 ;
  assign n16520 = n16443 & n16519 ;
  assign n16521 = n16520 ^ n14520 ;
  assign n16616 = n16521 ^ n14582 ;
  assign n16424 = n16082 ^ n16080 ;
  assign n16419 = n16418 ^ n15624 ;
  assign n16420 = ~n16417 & n16419 ;
  assign n16405 = n15624 ^ n15619 ;
  assign n16421 = n16420 ^ n16405 ;
  assign n16434 = n16424 ^ n16421 ;
  assign n16435 = n16434 ^ n15619 ;
  assign n16436 = n15280 & ~n16435 ;
  assign n16437 = n16436 ^ n15619 ;
  assign n16617 = n16616 ^ n16437 ;
  assign n16619 = n16617 ^ x467 ;
  assign n16618 = n16617 ^ n16610 ;
  assign n16620 = n16619 ^ n16618 ;
  assign n16621 = ~n16615 & n16620 ;
  assign n16622 = n16621 ^ n16619 ;
  assign n16438 = n16437 ^ n14582 ;
  assign n16522 = n16521 ^ n16437 ;
  assign n16523 = ~n16438 & ~n16522 ;
  assign n16524 = n16523 ^ n14582 ;
  assign n16623 = n16524 ^ n14628 ;
  assign n16428 = n16084 ^ n16083 ;
  assign n16422 = n15761 ^ n15619 ;
  assign n16423 = n16422 ^ n15761 ;
  assign n16425 = n16424 ^ n16423 ;
  assign n16426 = n16421 & ~n16425 ;
  assign n16427 = n16426 ^ n16422 ;
  assign n16429 = n16428 ^ n16427 ;
  assign n16430 = n16429 ^ n15761 ;
  assign n16431 = n15227 & ~n16430 ;
  assign n16432 = n16431 ^ n15761 ;
  assign n16624 = n16623 ^ n16432 ;
  assign n16626 = n16624 ^ x466 ;
  assign n16625 = n16624 ^ n16617 ;
  assign n16627 = n16626 ^ n16625 ;
  assign n16628 = ~n16622 & n16627 ;
  assign n16629 = n16628 ^ n16626 ;
  assign n16535 = n16086 ^ n16085 ;
  assign n16529 = n15912 ^ n15615 ;
  assign n16531 = n16529 ^ n15761 ;
  assign n16530 = n16529 ^ n16428 ;
  assign n16532 = n16531 ^ n16530 ;
  assign n16533 = n16427 & ~n16532 ;
  assign n16534 = n16533 ^ n16531 ;
  assign n16536 = n16535 ^ n16534 ;
  assign n16537 = n16536 ^ n16529 ;
  assign n16538 = n15295 & n16537 ;
  assign n16539 = n16538 ^ n16529 ;
  assign n16433 = n16432 ^ n14628 ;
  assign n16525 = n16524 ^ n16432 ;
  assign n16526 = n16433 & n16525 ;
  assign n16527 = n16526 ^ n14628 ;
  assign n16528 = n16527 ^ n14709 ;
  assign n16540 = n16539 ^ n16528 ;
  assign n16631 = n16540 ^ x465 ;
  assign n16630 = n16624 ^ n16540 ;
  assign n16632 = n16631 ^ n16630 ;
  assign n16633 = ~n16629 & n16632 ;
  assign n16634 = n16633 ^ n16631 ;
  assign n16810 = n16634 ^ x464 ;
  assign n16317 = n16316 ^ x462 ;
  assign n16318 = n16207 ^ x454 ;
  assign n16319 = n16318 ^ n16205 ;
  assign n16320 = n16221 ^ x453 ;
  assign n16321 = n16319 & n16320 ;
  assign n16322 = n16233 ^ x452 ;
  assign n16323 = ~n16321 & ~n16322 ;
  assign n16324 = n16245 ^ x451 ;
  assign n16325 = ~n16323 & n16324 ;
  assign n16326 = n16259 ^ x450 ;
  assign n16327 = ~n16325 & n16326 ;
  assign n16328 = n16272 ^ x449 ;
  assign n16329 = ~n16327 & ~n16328 ;
  assign n16330 = n16287 ^ x448 ;
  assign n16331 = n16329 & ~n16330 ;
  assign n16332 = n16302 ^ x463 ;
  assign n16333 = n16331 & ~n16332 ;
  assign n16782 = ~n16317 & n16333 ;
  assign n16783 = n16551 ^ x461 ;
  assign n16784 = n16782 & n16783 ;
  assign n16785 = n16558 ^ x460 ;
  assign n16786 = ~n16784 & n16785 ;
  assign n16787 = n16565 ^ x459 ;
  assign n16788 = n16786 & ~n16787 ;
  assign n16789 = n16572 ^ x458 ;
  assign n16790 = n16788 & ~n16789 ;
  assign n16791 = n16579 ^ x457 ;
  assign n16792 = n16790 & ~n16791 ;
  assign n16793 = n16584 ^ x456 ;
  assign n16794 = n16792 & n16793 ;
  assign n16795 = n16586 ^ x471 ;
  assign n16796 = n16795 ^ n16587 ;
  assign n16797 = ~n16794 & ~n16796 ;
  assign n16798 = n16594 ^ x470 ;
  assign n16799 = n16797 & ~n16798 ;
  assign n16800 = n16601 ^ x469 ;
  assign n16801 = n16799 & n16800 ;
  assign n16802 = n16608 ^ x468 ;
  assign n16803 = ~n16801 & n16802 ;
  assign n16804 = n16615 ^ x467 ;
  assign n16805 = ~n16803 & ~n16804 ;
  assign n16806 = n16622 ^ x466 ;
  assign n16807 = n16805 & ~n16806 ;
  assign n16808 = n16629 ^ x465 ;
  assign n16809 = ~n16807 & n16808 ;
  assign n16864 = n16810 ^ n16809 ;
  assign n16964 = ~n16142 & n16864 ;
  assign n16965 = n16964 ^ n16143 ;
  assign n17150 = n16965 ^ n15148 ;
  assign n17151 = x103 & n17150 ;
  assign n17355 = n17151 ^ x102 ;
  assign n16541 = n16540 ^ x464 ;
  assign n16635 = ~n16541 & n16634 ;
  assign n16636 = n16635 ^ x464 ;
  assign n16812 = n16636 ^ x479 ;
  assign n16637 = n16539 ^ n16527 ;
  assign n16644 = n16088 ^ n16087 ;
  assign n16638 = n15925 ^ n15915 ;
  assign n16640 = n16638 ^ n16529 ;
  assign n16639 = n16638 ^ n16535 ;
  assign n16641 = n16640 ^ n16639 ;
  assign n16642 = ~n16534 & ~n16641 ;
  assign n16643 = n16642 ^ n16640 ;
  assign n16645 = n16644 ^ n16643 ;
  assign n16646 = n16645 ^ n16638 ;
  assign n16647 = ~n15919 & n16646 ;
  assign n16648 = n16647 ^ n16638 ;
  assign n16649 = n16648 ^ n14709 ;
  assign n16650 = n16649 ^ n16527 ;
  assign n16651 = n16650 ^ n16648 ;
  assign n16652 = n16637 & ~n16651 ;
  assign n16653 = n16652 ^ n16649 ;
  assign n16654 = n16653 ^ n15230 ;
  assign n16813 = n16812 ^ n16654 ;
  assign n16811 = n16809 & ~n16810 ;
  assign n16868 = n16813 ^ n16811 ;
  assign n16863 = n16143 ^ n16142 ;
  assign n16865 = ~n16863 & ~n16864 ;
  assign n16869 = n16868 ^ n16865 ;
  assign n16968 = ~n16145 & ~n16869 ;
  assign n16866 = n16147 ^ n16146 ;
  assign n16969 = n16968 ^ n16866 ;
  assign n16966 = n15148 & n16965 ;
  assign n16967 = n16966 ^ n15152 ;
  assign n17149 = n16969 ^ n16967 ;
  assign n17356 = n17355 ^ n17149 ;
  assign n17354 = n17150 ^ x103 ;
  assign n17763 = n17356 ^ n17354 ;
  assign n16922 = n16328 ^ n16327 ;
  assign n16898 = n16307 ^ n16196 ;
  assign n16893 = n16307 ^ n16288 ;
  assign n16655 = n16654 ^ n16636 ;
  assign n16657 = n16644 ^ n16638 ;
  assign n16658 = ~n16643 & ~n16657 ;
  assign n16659 = n16658 ^ n16638 ;
  assign n16656 = n16090 ^ n16089 ;
  assign n16660 = n16659 ^ n16656 ;
  assign n16661 = ~n15943 & ~n16660 ;
  assign n16662 = n16661 ^ n15929 ;
  assign n16664 = n16662 ^ n15230 ;
  assign n16663 = n16662 ^ n16648 ;
  assign n16665 = n16664 ^ n16663 ;
  assign n16666 = n16653 & n16665 ;
  assign n16667 = n16666 ^ n16664 ;
  assign n16668 = n16667 ^ n15310 ;
  assign n16669 = n16668 ^ x479 ;
  assign n16670 = n16669 ^ n16636 ;
  assign n16671 = n16670 ^ n16668 ;
  assign n16672 = ~n16655 & n16671 ;
  assign n16673 = n16672 ^ n16669 ;
  assign n16683 = n16092 ^ n16091 ;
  assign n16681 = n16656 ^ n15952 ;
  assign n16678 = n15943 ^ n15929 ;
  assign n16679 = n16678 ^ n16656 ;
  assign n16680 = n16660 & n16679 ;
  assign n16682 = n16681 ^ n16680 ;
  assign n16684 = n16683 ^ n16682 ;
  assign n16685 = n16684 ^ n15952 ;
  assign n16686 = ~n15945 & ~n16685 ;
  assign n16687 = n16686 ^ n15952 ;
  assign n16674 = n16662 ^ n15310 ;
  assign n16675 = n16667 & n16674 ;
  assign n16676 = n16675 ^ n15310 ;
  assign n16677 = n16676 ^ n15325 ;
  assign n16688 = n16687 ^ n16677 ;
  assign n16690 = n16688 ^ x478 ;
  assign n16689 = n16688 ^ n16668 ;
  assign n16691 = n16690 ^ n16689 ;
  assign n16692 = n16673 & ~n16691 ;
  assign n16693 = n16692 ^ n16690 ;
  assign n16704 = n16094 ^ n16093 ;
  assign n16700 = n15976 ^ n15952 ;
  assign n16699 = n16683 ^ n15976 ;
  assign n16701 = n16700 ^ n16699 ;
  assign n16702 = ~n16682 & n16701 ;
  assign n16703 = n16702 ^ n16700 ;
  assign n16705 = n16704 ^ n16703 ;
  assign n16706 = n16705 ^ n15976 ;
  assign n16707 = n15330 & n16706 ;
  assign n16708 = n16707 ^ n15976 ;
  assign n16694 = n16687 ^ n16676 ;
  assign n16695 = n16687 ^ n15325 ;
  assign n16696 = ~n16694 & n16695 ;
  assign n16697 = n16696 ^ n15325 ;
  assign n16698 = n16697 ^ n14873 ;
  assign n16709 = n16708 ^ n16698 ;
  assign n16711 = n16709 ^ x477 ;
  assign n16710 = n16709 ^ n16688 ;
  assign n16712 = n16711 ^ n16710 ;
  assign n16713 = ~n16693 & n16712 ;
  assign n16714 = n16713 ^ n16711 ;
  assign n16725 = n16096 ^ n16095 ;
  assign n16721 = n15997 ^ n15976 ;
  assign n16720 = n16704 ^ n15997 ;
  assign n16722 = n16721 ^ n16720 ;
  assign n16723 = n16703 & n16722 ;
  assign n16724 = n16723 ^ n16721 ;
  assign n16726 = n16725 ^ n16724 ;
  assign n16727 = n16726 ^ n15997 ;
  assign n16728 = n15344 & ~n16727 ;
  assign n16729 = n16728 ^ n15997 ;
  assign n16715 = n16708 ^ n16697 ;
  assign n16716 = n16708 ^ n14873 ;
  assign n16717 = ~n16715 & n16716 ;
  assign n16718 = n16717 ^ n14873 ;
  assign n16719 = n16718 ^ n14914 ;
  assign n16730 = n16729 ^ n16719 ;
  assign n16732 = n16730 ^ x476 ;
  assign n16731 = n16730 ^ n16709 ;
  assign n16733 = n16732 ^ n16731 ;
  assign n16734 = ~n16714 & n16733 ;
  assign n16735 = n16734 ^ n16732 ;
  assign n16746 = n16099 ^ n16097 ;
  assign n16742 = n16018 ^ n15997 ;
  assign n16741 = n16725 ^ n16018 ;
  assign n16743 = n16742 ^ n16741 ;
  assign n16744 = n16724 & ~n16743 ;
  assign n16745 = n16744 ^ n16742 ;
  assign n16747 = n16746 ^ n16745 ;
  assign n16748 = n16747 ^ n16018 ;
  assign n16749 = n15358 & ~n16748 ;
  assign n16750 = n16749 ^ n16018 ;
  assign n16736 = n16729 ^ n16718 ;
  assign n16737 = n16729 ^ n14914 ;
  assign n16738 = ~n16736 & ~n16737 ;
  assign n16739 = n16738 ^ n14914 ;
  assign n16740 = n16739 ^ n14954 ;
  assign n16751 = n16750 ^ n16740 ;
  assign n16753 = n16751 ^ x475 ;
  assign n16752 = n16751 ^ n16730 ;
  assign n16754 = n16753 ^ n16752 ;
  assign n16755 = n16735 & ~n16754 ;
  assign n16756 = n16755 ^ n16753 ;
  assign n16767 = n16101 ^ n16100 ;
  assign n16763 = n16039 ^ n16018 ;
  assign n16762 = n16746 ^ n16039 ;
  assign n16764 = n16763 ^ n16762 ;
  assign n16765 = n16745 & ~n16764 ;
  assign n16766 = n16765 ^ n16763 ;
  assign n16768 = n16767 ^ n16766 ;
  assign n16769 = n16768 ^ n16039 ;
  assign n16770 = ~n15372 & n16769 ;
  assign n16771 = n16770 ^ n16039 ;
  assign n16757 = n16750 ^ n16739 ;
  assign n16758 = n16750 ^ n14954 ;
  assign n16759 = n16757 & n16758 ;
  assign n16760 = n16759 ^ n14954 ;
  assign n16761 = n16760 ^ n14990 ;
  assign n16772 = n16771 ^ n16761 ;
  assign n16774 = n16772 ^ x474 ;
  assign n16773 = n16772 ^ n16751 ;
  assign n16775 = n16774 ^ n16773 ;
  assign n16776 = n16756 & ~n16775 ;
  assign n16777 = n16776 ^ n16774 ;
  assign n16844 = n16777 ^ x473 ;
  assign n16779 = n16735 ^ x475 ;
  assign n16780 = n16714 ^ x476 ;
  assign n16781 = n16693 ^ x477 ;
  assign n16814 = ~n16811 & ~n16813 ;
  assign n16815 = n16673 ^ x478 ;
  assign n16816 = n16814 & n16815 ;
  assign n16817 = n16781 & ~n16816 ;
  assign n16818 = n16780 & n16817 ;
  assign n16819 = ~n16779 & n16818 ;
  assign n16820 = n16756 ^ x474 ;
  assign n16821 = n16819 & ~n16820 ;
  assign n16845 = n16844 ^ n16821 ;
  assign n16846 = n16845 ^ n16278 ;
  assign n16848 = n16165 ^ n16052 ;
  assign n16847 = n16820 ^ n16819 ;
  assign n16849 = n16848 ^ n16847 ;
  assign n16850 = n16818 ^ n16779 ;
  assign n16851 = n16850 ^ n16246 ;
  assign n16854 = n16817 ^ n16780 ;
  assign n16852 = n16156 ^ n16132 ;
  assign n16853 = n16852 ^ n16131 ;
  assign n16855 = n16854 ^ n16853 ;
  assign n16857 = n16153 ^ n16137 ;
  assign n16858 = n16857 ^ n16135 ;
  assign n16856 = n16816 ^ n16781 ;
  assign n16859 = n16858 ^ n16856 ;
  assign n16861 = n16815 ^ n16814 ;
  assign n16860 = n16151 ^ n16140 ;
  assign n16862 = n16861 ^ n16860 ;
  assign n16867 = n16866 ^ n16865 ;
  assign n16870 = n16867 & n16869 ;
  assign n16871 = n16870 ^ n16866 ;
  assign n16872 = n16871 ^ n16860 ;
  assign n16873 = n16862 & n16872 ;
  assign n16874 = n16873 ^ n16861 ;
  assign n16875 = n16874 ^ n16856 ;
  assign n16876 = n16859 & ~n16875 ;
  assign n16877 = n16876 ^ n16858 ;
  assign n16878 = n16877 ^ n16853 ;
  assign n16879 = ~n16855 & ~n16878 ;
  assign n16880 = n16879 ^ n16854 ;
  assign n16881 = n16880 ^ n16850 ;
  assign n16882 = ~n16851 & n16881 ;
  assign n16883 = n16882 ^ n16246 ;
  assign n16884 = n16883 ^ n16847 ;
  assign n16885 = ~n16849 & n16884 ;
  assign n16886 = n16885 ^ n16848 ;
  assign n16887 = n16886 ^ n16845 ;
  assign n16888 = n16846 & ~n16887 ;
  assign n16889 = n16888 ^ n16278 ;
  assign n16837 = n16767 ^ n16039 ;
  assign n16838 = ~n16766 & n16837 ;
  assign n16835 = n16103 ^ n16102 ;
  assign n16834 = n16767 ^ n16127 ;
  assign n16836 = n16835 ^ n16834 ;
  assign n16839 = n16838 ^ n16836 ;
  assign n16840 = n16839 ^ n16127 ;
  assign n16841 = n15388 & n16840 ;
  assign n16831 = n16127 ^ n15041 ;
  assign n16830 = n14990 ^ x472 ;
  assign n16832 = n16831 ^ n16830 ;
  assign n16827 = n16771 ^ n16760 ;
  assign n16828 = n16771 ^ n14990 ;
  assign n16829 = ~n16827 & ~n16828 ;
  assign n16833 = n16832 ^ n16829 ;
  assign n16842 = n16841 ^ n16833 ;
  assign n16822 = n16821 ^ n16772 ;
  assign n16825 = n16777 & n16822 ;
  assign n16778 = n16777 ^ n16772 ;
  assign n16823 = n16822 ^ n16778 ;
  assign n16824 = x473 & n16823 ;
  assign n16826 = n16825 ^ n16824 ;
  assign n16843 = n16842 ^ n16826 ;
  assign n16890 = n16889 ^ n16843 ;
  assign n16891 = n16889 ^ n16288 ;
  assign n16892 = ~n16890 & n16891 ;
  assign n16894 = n16893 ^ n16892 ;
  assign n16895 = n16206 ^ x455 ;
  assign n16896 = n16895 ^ n16307 ;
  assign n16897 = n16894 & ~n16896 ;
  assign n16899 = n16898 ^ n16897 ;
  assign n16900 = n16319 ^ n16196 ;
  assign n16901 = ~n16899 & ~n16900 ;
  assign n16404 = n16402 ^ n16196 ;
  assign n16902 = n16901 ^ n16404 ;
  assign n16903 = n16320 ^ n16319 ;
  assign n16904 = n16903 ^ n16402 ;
  assign n16905 = n16902 & n16904 ;
  assign n16403 = n16402 ^ n16400 ;
  assign n16906 = n16905 ^ n16403 ;
  assign n16907 = n16322 ^ n16321 ;
  assign n16908 = n16907 ^ n16400 ;
  assign n16909 = n16906 & ~n16908 ;
  assign n16401 = n16400 ^ n16398 ;
  assign n16910 = n16909 ^ n16401 ;
  assign n16911 = n16324 ^ n16323 ;
  assign n16912 = n16911 ^ n16398 ;
  assign n16913 = ~n16910 & n16912 ;
  assign n16399 = n16398 ^ n16395 ;
  assign n16914 = n16913 ^ n16399 ;
  assign n16915 = n16326 ^ n16325 ;
  assign n16916 = n16915 ^ n16395 ;
  assign n16917 = n16914 & ~n16916 ;
  assign n16397 = n16396 ^ n16395 ;
  assign n16918 = n16917 ^ n16397 ;
  assign n17042 = n16922 ^ n16918 ;
  assign n16939 = n16915 ^ n16914 ;
  assign n17761 = n17042 ^ n16939 ;
  assign n17127 = n16536 ^ n16429 ;
  assign n16393 = n16332 ^ n16331 ;
  assign n16385 = n16384 ^ n16383 ;
  assign n16394 = n16393 ^ n16385 ;
  assign n16919 = n16378 ^ n16377 ;
  assign n16920 = n16919 ^ n16396 ;
  assign n16921 = n16920 ^ n16919 ;
  assign n16923 = n16922 ^ n16921 ;
  assign n16924 = n16918 & ~n16923 ;
  assign n16925 = n16924 ^ n16920 ;
  assign n16928 = n16919 ^ n16385 ;
  assign n16926 = n16330 ^ n16329 ;
  assign n16927 = n16926 ^ n16385 ;
  assign n16929 = n16928 ^ n16927 ;
  assign n16930 = n16925 & n16929 ;
  assign n16931 = n16930 ^ n16928 ;
  assign n16932 = ~n16394 & ~n16931 ;
  assign n16392 = n16391 ^ n16385 ;
  assign n16933 = n16932 ^ n16392 ;
  assign n16334 = n16333 ^ n16317 ;
  assign n17074 = n16391 ^ n16334 ;
  assign n17075 = n16933 & ~n17074 ;
  assign n17073 = n16444 ^ n16391 ;
  assign n17076 = n17075 ^ n17073 ;
  assign n17072 = n16783 ^ n16782 ;
  assign n17087 = n17072 ^ n16444 ;
  assign n17088 = ~n17076 & ~n17087 ;
  assign n17086 = n16444 ^ n16439 ;
  assign n17089 = n17088 ^ n17086 ;
  assign n17085 = n16785 ^ n16784 ;
  assign n17100 = n17085 ^ n16439 ;
  assign n17101 = n17089 & ~n17100 ;
  assign n17099 = n16439 ^ n16434 ;
  assign n17102 = n17101 ^ n17099 ;
  assign n17098 = n16787 ^ n16786 ;
  assign n17113 = n17098 ^ n16434 ;
  assign n17114 = n17102 & ~n17113 ;
  assign n17112 = n16434 ^ n16429 ;
  assign n17115 = n17114 ^ n17112 ;
  assign n17111 = n16789 ^ n16788 ;
  assign n17125 = n17111 ^ n16429 ;
  assign n17126 = n17115 & ~n17125 ;
  assign n17128 = n17127 ^ n17126 ;
  assign n17124 = n16791 ^ n16790 ;
  assign n17129 = n17128 ^ n17124 ;
  assign n17130 = n17129 ^ n16536 ;
  assign n17131 = n16529 & ~n17130 ;
  assign n17132 = n17131 ^ n16536 ;
  assign n16934 = n16933 ^ n16334 ;
  assign n16935 = n16934 ^ n16391 ;
  assign n16936 = n16198 & ~n16935 ;
  assign n16937 = n16936 ^ n16391 ;
  assign n16938 = n16937 ^ n15252 ;
  assign n17059 = n16931 ^ n16393 ;
  assign n17060 = n17059 ^ n16383 ;
  assign n17061 = ~n16384 & n17060 ;
  assign n17062 = n17061 ^ n17059 ;
  assign n17043 = n17042 ^ n16396 ;
  assign n17044 = ~n16366 & ~n17043 ;
  assign n17045 = n17044 ^ n16396 ;
  assign n16940 = n16939 ^ n16395 ;
  assign n16941 = ~n16358 & ~n16940 ;
  assign n16942 = n16941 ^ n16395 ;
  assign n16943 = n16942 ^ n15516 ;
  assign n16944 = n16911 ^ n16910 ;
  assign n16945 = n16944 ^ n16398 ;
  assign n16946 = ~n16351 & ~n16945 ;
  assign n16947 = n16946 ^ n16398 ;
  assign n16948 = n16947 ^ n15521 ;
  assign n16949 = n16907 ^ n16906 ;
  assign n16950 = n16949 ^ n16400 ;
  assign n16951 = n16343 & ~n16950 ;
  assign n16952 = n16951 ^ n16400 ;
  assign n16953 = n16952 ^ n15524 ;
  assign n16954 = n16903 ^ n16902 ;
  assign n16955 = n16954 ^ n16402 ;
  assign n16956 = n16336 & n16955 ;
  assign n16957 = n16956 ^ n16402 ;
  assign n16958 = n16957 ^ n15529 ;
  assign n17022 = n16899 ^ n16319 ;
  assign n17023 = n17022 ^ n16196 ;
  assign n17024 = n16189 & n17023 ;
  assign n17025 = n17024 ^ n16196 ;
  assign n16959 = n15191 & ~n16881 ;
  assign n16960 = n16959 ^ n16246 ;
  assign n16961 = n16960 ^ n15168 ;
  assign n16970 = n16969 ^ n16966 ;
  assign n16971 = ~n16967 & ~n16970 ;
  assign n16972 = n16971 ^ n15152 ;
  assign n16973 = n16972 ^ n15145 ;
  assign n16974 = n16871 ^ n16861 ;
  assign n16975 = ~n16139 & ~n16974 ;
  assign n16976 = n16975 ^ n16860 ;
  assign n16977 = n16976 ^ n16972 ;
  assign n16978 = n16973 & ~n16977 ;
  assign n16979 = n16978 ^ n15145 ;
  assign n16962 = n16137 & n16875 ;
  assign n16963 = n16962 ^ n16858 ;
  assign n16980 = n16979 ^ n16963 ;
  assign n16981 = n16877 ^ n16854 ;
  assign n16982 = n16132 & ~n16981 ;
  assign n16983 = n16982 ^ n16853 ;
  assign n16984 = n16983 ^ n15142 ;
  assign n16985 = n16984 ^ n16963 ;
  assign n16986 = n16985 ^ n16983 ;
  assign n16987 = ~n16980 & ~n16986 ;
  assign n16988 = n16987 ^ n16984 ;
  assign n16990 = n16960 ^ n14644 ;
  assign n16989 = n16983 ^ n16960 ;
  assign n16991 = n16990 ^ n16989 ;
  assign n16992 = n16988 & ~n16991 ;
  assign n16993 = n16992 ^ n16990 ;
  assign n16994 = n16961 & ~n16993 ;
  assign n16995 = n16994 ^ n15168 ;
  assign n16996 = n16995 ^ n15549 ;
  assign n16997 = ~n16164 & ~n16884 ;
  assign n16998 = n16997 ^ n16848 ;
  assign n16999 = n16998 ^ n16995 ;
  assign n17000 = n16996 & ~n16999 ;
  assign n17001 = n17000 ^ n15549 ;
  assign n17002 = n17001 ^ n15545 ;
  assign n17003 = n16167 & n16887 ;
  assign n17004 = n17003 ^ n16278 ;
  assign n17005 = n17004 ^ n17001 ;
  assign n17006 = n17002 & ~n17005 ;
  assign n17007 = n17006 ^ n15545 ;
  assign n17008 = n17007 ^ n15540 ;
  assign n17009 = n16174 & n16890 ;
  assign n17010 = n17009 ^ n16288 ;
  assign n17011 = n17010 ^ n17007 ;
  assign n17012 = ~n17008 & ~n17011 ;
  assign n17013 = n17012 ^ n15540 ;
  assign n17014 = n17013 ^ n15537 ;
  assign n17015 = n16895 ^ n16894 ;
  assign n17016 = n17015 ^ n16307 ;
  assign n17017 = ~n16182 & ~n17016 ;
  assign n17018 = n17017 ^ n16307 ;
  assign n17019 = n17018 ^ n17013 ;
  assign n17020 = n17014 & n17019 ;
  assign n17021 = n17020 ^ n15537 ;
  assign n17026 = n17025 ^ n17021 ;
  assign n17027 = n17025 ^ n15532 ;
  assign n17028 = ~n17026 & n17027 ;
  assign n17029 = n17028 ^ n15532 ;
  assign n17030 = n17029 ^ n16957 ;
  assign n17031 = ~n16958 & ~n17030 ;
  assign n17032 = n17031 ^ n15529 ;
  assign n17033 = n17032 ^ n16952 ;
  assign n17034 = n16953 & n17033 ;
  assign n17035 = n17034 ^ n15524 ;
  assign n17036 = n17035 ^ n16947 ;
  assign n17037 = ~n16948 & n17036 ;
  assign n17038 = n17037 ^ n15521 ;
  assign n17039 = n17038 ^ n16942 ;
  assign n17040 = ~n16943 & n17039 ;
  assign n17041 = n17040 ^ n15516 ;
  assign n17046 = n17045 ^ n17041 ;
  assign n17047 = n16926 ^ n16925 ;
  assign n17048 = n17047 ^ n16377 ;
  assign n17049 = n16378 & n17048 ;
  assign n17050 = n17049 ^ n16377 ;
  assign n17051 = n17050 ^ n15083 ;
  assign n17052 = n17051 ^ n17041 ;
  assign n17053 = n17052 ^ n17050 ;
  assign n17054 = n17046 & n17053 ;
  assign n17055 = n17054 ^ n17051 ;
  assign n17056 = n17050 ^ n15586 ;
  assign n17057 = n17055 & n17056 ;
  assign n17058 = n17057 ^ n15586 ;
  assign n17063 = n17062 ^ n17058 ;
  assign n17064 = n16937 ^ n15512 ;
  assign n17065 = n17064 ^ n17058 ;
  assign n17066 = n17065 ^ n16937 ;
  assign n17067 = n17063 & ~n17066 ;
  assign n17068 = n17067 ^ n17064 ;
  assign n17069 = ~n16938 & ~n17068 ;
  assign n17070 = n17069 ^ n15252 ;
  assign n17071 = n17070 ^ n15507 ;
  assign n17077 = n17076 ^ n17072 ;
  assign n17078 = n17077 ^ n16444 ;
  assign n17079 = n16407 & n17078 ;
  assign n17080 = n17079 ^ n16444 ;
  assign n17081 = n17080 ^ n17070 ;
  assign n17082 = ~n17071 & ~n17081 ;
  assign n17083 = n17082 ^ n15507 ;
  assign n17084 = n17083 ^ n15272 ;
  assign n17090 = n17089 ^ n17085 ;
  assign n17091 = n17090 ^ n16439 ;
  assign n17092 = ~n15624 & ~n17091 ;
  assign n17093 = n17092 ^ n16439 ;
  assign n17094 = n17093 ^ n17083 ;
  assign n17095 = ~n17084 & n17094 ;
  assign n17096 = n17095 ^ n15272 ;
  assign n17097 = n17096 ^ n15280 ;
  assign n17103 = n17102 ^ n17098 ;
  assign n17104 = n17103 ^ n16434 ;
  assign n17105 = ~n15619 & ~n17104 ;
  assign n17106 = n17105 ^ n16434 ;
  assign n17107 = n17106 ^ n17096 ;
  assign n17108 = n17097 & ~n17107 ;
  assign n17109 = n17108 ^ n15280 ;
  assign n17110 = n17109 ^ n15227 ;
  assign n17116 = n17115 ^ n17111 ;
  assign n17117 = n17116 ^ n16429 ;
  assign n17118 = ~n15761 & ~n17117 ;
  assign n17119 = n17118 ^ n16429 ;
  assign n17120 = n17119 ^ n17109 ;
  assign n17121 = n17110 & ~n17120 ;
  assign n17122 = n17121 ^ n15227 ;
  assign n17276 = n17132 ^ n17122 ;
  assign n17277 = n16793 ^ n16792 ;
  assign n17278 = n17277 ^ n16536 ;
  assign n17279 = n17278 ^ n17124 ;
  assign n17280 = n17279 ^ n17277 ;
  assign n17281 = n17128 & ~n17280 ;
  assign n17282 = n17281 ^ n17278 ;
  assign n17283 = ~n16638 & n17282 ;
  assign n17284 = n17283 ^ n16645 ;
  assign n17285 = n17284 ^ n15295 ;
  assign n17286 = n17285 ^ n17122 ;
  assign n17287 = n17286 ^ n17284 ;
  assign n17288 = ~n17276 & n17287 ;
  assign n17289 = n17288 ^ n17285 ;
  assign n17290 = n17289 ^ n15919 ;
  assign n17123 = n17122 ^ n15295 ;
  assign n17133 = n17132 ^ n17123 ;
  assign n17134 = n17133 ^ x112 ;
  assign n17243 = n17068 ^ n15252 ;
  assign n17135 = n17058 ^ n15512 ;
  assign n17136 = n17135 ^ n17062 ;
  assign n17137 = n17136 ^ x118 ;
  assign n17234 = n17055 ^ n15586 ;
  assign n17138 = n17041 ^ n15083 ;
  assign n17139 = n17138 ^ n17045 ;
  assign n17140 = n17139 ^ x104 ;
  assign n17141 = n17038 ^ n15516 ;
  assign n17142 = n17141 ^ n16942 ;
  assign n17143 = n17142 ^ x105 ;
  assign n17146 = n17021 ^ n15532 ;
  assign n17147 = n17146 ^ n17025 ;
  assign n17148 = n17147 ^ x109 ;
  assign n17152 = n17151 ^ n17149 ;
  assign n17153 = n16976 ^ n16973 ;
  assign n17154 = n17153 ^ x102 ;
  assign n17155 = n17154 ^ n17149 ;
  assign n17156 = n17155 ^ n17153 ;
  assign n17157 = n17152 & ~n17156 ;
  assign n17158 = n17157 ^ n17154 ;
  assign n17159 = n16979 ^ n15142 ;
  assign n17160 = n17159 ^ n16963 ;
  assign n17162 = n17160 ^ x101 ;
  assign n17161 = n17160 ^ n17153 ;
  assign n17163 = n17162 ^ n17161 ;
  assign n17164 = n17158 & ~n17163 ;
  assign n17165 = n17164 ^ n17162 ;
  assign n17166 = n16988 ^ n14644 ;
  assign n17168 = n17166 ^ x100 ;
  assign n17167 = n17166 ^ n17160 ;
  assign n17169 = n17168 ^ n17167 ;
  assign n17170 = ~n17165 & n17169 ;
  assign n17171 = n17170 ^ n17168 ;
  assign n17172 = n16993 ^ n15168 ;
  assign n17174 = n17172 ^ x99 ;
  assign n17173 = n17172 ^ n17166 ;
  assign n17175 = n17174 ^ n17173 ;
  assign n17176 = n17171 & ~n17175 ;
  assign n17177 = n17176 ^ n17174 ;
  assign n17178 = n16998 ^ n16996 ;
  assign n17180 = n17178 ^ x98 ;
  assign n17179 = n17178 ^ n17172 ;
  assign n17181 = n17180 ^ n17179 ;
  assign n17182 = ~n17177 & n17181 ;
  assign n17183 = n17182 ^ n17180 ;
  assign n17184 = n17004 ^ n17002 ;
  assign n17186 = n17184 ^ x97 ;
  assign n17185 = n17184 ^ n17178 ;
  assign n17187 = n17186 ^ n17185 ;
  assign n17188 = ~n17183 & n17187 ;
  assign n17189 = n17188 ^ n17186 ;
  assign n17190 = n17010 ^ n17008 ;
  assign n17192 = n17190 ^ x96 ;
  assign n17191 = n17190 ^ n17184 ;
  assign n17193 = n17192 ^ n17191 ;
  assign n17194 = ~n17189 & n17193 ;
  assign n17195 = n17194 ^ n17192 ;
  assign n17196 = n17018 ^ n17014 ;
  assign n17198 = n17196 ^ x111 ;
  assign n17197 = n17196 ^ n17190 ;
  assign n17199 = n17198 ^ n17197 ;
  assign n17200 = n17195 & ~n17199 ;
  assign n17201 = n17200 ^ n17198 ;
  assign n17203 = n17147 ^ x110 ;
  assign n17202 = n17196 ^ n17147 ;
  assign n17204 = n17203 ^ n17202 ;
  assign n17205 = ~n17201 & n17204 ;
  assign n17206 = n17205 ^ n17203 ;
  assign n17207 = ~n17148 & n17206 ;
  assign n17208 = n17207 ^ x109 ;
  assign n17144 = n17029 ^ n15529 ;
  assign n17145 = n17144 ^ n16957 ;
  assign n17209 = n17208 ^ n17145 ;
  assign n17210 = n17032 ^ n15524 ;
  assign n17211 = n17210 ^ n16952 ;
  assign n17212 = n17211 ^ x108 ;
  assign n17213 = n17212 ^ n17208 ;
  assign n17214 = n17213 ^ n17211 ;
  assign n17215 = ~n17209 & n17214 ;
  assign n17216 = n17215 ^ n17212 ;
  assign n17217 = n17035 ^ n15521 ;
  assign n17218 = n17217 ^ n16947 ;
  assign n17220 = n17218 ^ x107 ;
  assign n17219 = n17218 ^ n17211 ;
  assign n17221 = n17220 ^ n17219 ;
  assign n17222 = ~n17216 & n17221 ;
  assign n17223 = n17222 ^ n17220 ;
  assign n17225 = n17142 ^ x106 ;
  assign n17224 = n17218 ^ n17142 ;
  assign n17226 = n17225 ^ n17224 ;
  assign n17227 = ~n17223 & n17226 ;
  assign n17228 = n17227 ^ n17225 ;
  assign n17229 = n17143 & ~n17228 ;
  assign n17230 = n17229 ^ x105 ;
  assign n17231 = n17230 ^ n17139 ;
  assign n17232 = n17140 & ~n17231 ;
  assign n17233 = n17232 ^ x104 ;
  assign n17235 = n17234 ^ n17233 ;
  assign n17236 = n17136 ^ x119 ;
  assign n17237 = n17236 ^ n17136 ;
  assign n17238 = n17237 ^ n17233 ;
  assign n17239 = n17235 & n17238 ;
  assign n17240 = n17239 ^ n17236 ;
  assign n17241 = n17137 & ~n17240 ;
  assign n17242 = n17241 ^ x118 ;
  assign n17244 = n17243 ^ n17242 ;
  assign n17245 = n17080 ^ n17071 ;
  assign n17246 = n17245 ^ x117 ;
  assign n17247 = n17246 ^ n17242 ;
  assign n17248 = n17247 ^ n17245 ;
  assign n17249 = ~n17244 & n17248 ;
  assign n17250 = n17249 ^ n17246 ;
  assign n17251 = n17093 ^ n17084 ;
  assign n17253 = n17251 ^ x116 ;
  assign n17252 = n17251 ^ n17245 ;
  assign n17254 = n17253 ^ n17252 ;
  assign n17255 = n17250 & ~n17254 ;
  assign n17256 = n17255 ^ n17253 ;
  assign n17257 = n17106 ^ n17097 ;
  assign n17259 = n17257 ^ x115 ;
  assign n17258 = n17257 ^ n17251 ;
  assign n17260 = n17259 ^ n17258 ;
  assign n17261 = n17256 & ~n17260 ;
  assign n17262 = n17261 ^ n17259 ;
  assign n17263 = n17119 ^ n17110 ;
  assign n17265 = n17263 ^ x114 ;
  assign n17264 = n17263 ^ n17257 ;
  assign n17266 = n17265 ^ n17264 ;
  assign n17267 = ~n17262 & n17266 ;
  assign n17268 = n17267 ^ n17265 ;
  assign n17270 = n17133 ^ x113 ;
  assign n17269 = n17263 ^ n17133 ;
  assign n17271 = n17270 ^ n17269 ;
  assign n17272 = ~n17268 & n17271 ;
  assign n17273 = n17272 ^ n17270 ;
  assign n17274 = n17134 & ~n17273 ;
  assign n17275 = n17274 ^ x112 ;
  assign n17291 = n17290 ^ n17275 ;
  assign n17293 = n17277 ^ n16645 ;
  assign n17294 = ~n17282 & ~n17293 ;
  assign n17295 = n17294 ^ n16645 ;
  assign n17292 = n16796 ^ n16794 ;
  assign n17296 = n17295 ^ n17292 ;
  assign n17297 = ~n16678 & ~n17296 ;
  assign n17298 = n17297 ^ n16660 ;
  assign n17300 = n17298 ^ n15919 ;
  assign n17299 = n17298 ^ n17284 ;
  assign n17301 = n17300 ^ n17299 ;
  assign n17302 = n17289 & n17301 ;
  assign n17303 = n17302 ^ n17300 ;
  assign n17304 = n17303 ^ n15943 ;
  assign n17305 = n17304 ^ x127 ;
  assign n17306 = n17305 ^ n17275 ;
  assign n17307 = n17306 ^ n17304 ;
  assign n17308 = ~n17291 & n17307 ;
  assign n17309 = n17308 ^ n17305 ;
  assign n17319 = n16798 ^ n16797 ;
  assign n17317 = n17292 ^ n16684 ;
  assign n17314 = n16678 ^ n16660 ;
  assign n17315 = n17314 ^ n17292 ;
  assign n17316 = n17296 & n17315 ;
  assign n17318 = n17317 ^ n17316 ;
  assign n17320 = n17319 ^ n17318 ;
  assign n17321 = n17320 ^ n16684 ;
  assign n17322 = n15952 & ~n17321 ;
  assign n17323 = n17322 ^ n16684 ;
  assign n17310 = n17298 ^ n15943 ;
  assign n17311 = n17303 & ~n17310 ;
  assign n17312 = n17311 ^ n15943 ;
  assign n17313 = n17312 ^ n15945 ;
  assign n17324 = n17323 ^ n17313 ;
  assign n17326 = n17324 ^ x126 ;
  assign n17325 = n17324 ^ n17304 ;
  assign n17327 = n17326 ^ n17325 ;
  assign n17328 = ~n17309 & n17327 ;
  assign n17329 = n17328 ^ n17326 ;
  assign n17340 = n16800 ^ n16799 ;
  assign n17336 = n16705 ^ n16684 ;
  assign n17335 = n17319 ^ n16705 ;
  assign n17337 = n17336 ^ n17335 ;
  assign n17338 = n17318 & ~n17337 ;
  assign n17339 = n17338 ^ n17336 ;
  assign n17341 = n17340 ^ n17339 ;
  assign n17342 = n17341 ^ n16705 ;
  assign n17343 = n15976 & n17342 ;
  assign n17344 = n17343 ^ n16705 ;
  assign n17330 = n17323 ^ n17312 ;
  assign n17331 = n17323 ^ n15945 ;
  assign n17332 = ~n17330 & n17331 ;
  assign n17333 = n17332 ^ n15945 ;
  assign n17334 = n17333 ^ n15330 ;
  assign n17345 = n17344 ^ n17334 ;
  assign n17347 = n17345 ^ x125 ;
  assign n17346 = n17345 ^ n17324 ;
  assign n17348 = n17347 ^ n17346 ;
  assign n17349 = n17329 & ~n17348 ;
  assign n17350 = n17349 ^ n17347 ;
  assign n17479 = n16802 ^ n16801 ;
  assign n17475 = n16726 ^ n16705 ;
  assign n17474 = n17340 ^ n16726 ;
  assign n17476 = n17475 ^ n17474 ;
  assign n17477 = ~n17339 & ~n17476 ;
  assign n17478 = n17477 ^ n17475 ;
  assign n17480 = n17479 ^ n17478 ;
  assign n17481 = n17480 ^ n16726 ;
  assign n17482 = n15997 & ~n17481 ;
  assign n17483 = n17482 ^ n16726 ;
  assign n17469 = n17344 ^ n17333 ;
  assign n17470 = n17344 ^ n15330 ;
  assign n17471 = n17469 & n17470 ;
  assign n17472 = n17471 ^ n15330 ;
  assign n17473 = n17472 ^ n15344 ;
  assign n17484 = n17483 ^ n17473 ;
  assign n17486 = n17484 ^ x124 ;
  assign n17485 = n17484 ^ n17345 ;
  assign n17487 = n17486 ^ n17485 ;
  assign n17488 = n17350 & ~n17487 ;
  assign n17489 = n17488 ^ n17486 ;
  assign n17571 = n16804 ^ n16803 ;
  assign n17567 = n16747 ^ n16726 ;
  assign n17566 = n17479 ^ n16747 ;
  assign n17568 = n17567 ^ n17566 ;
  assign n17569 = ~n17478 & n17568 ;
  assign n17570 = n17569 ^ n17567 ;
  assign n17572 = n17571 ^ n17570 ;
  assign n17573 = n17572 ^ n16747 ;
  assign n17574 = n16018 & n17573 ;
  assign n17575 = n17574 ^ n16747 ;
  assign n17561 = n17483 ^ n17472 ;
  assign n17562 = n17483 ^ n15344 ;
  assign n17563 = n17561 & ~n17562 ;
  assign n17564 = n17563 ^ n15344 ;
  assign n17565 = n17564 ^ n15358 ;
  assign n17576 = n17575 ^ n17565 ;
  assign n17578 = n17576 ^ x123 ;
  assign n17577 = n17576 ^ n17484 ;
  assign n17579 = n17578 ^ n17577 ;
  assign n17580 = n17489 & ~n17579 ;
  assign n17581 = n17580 ^ n17578 ;
  assign n17683 = n16806 ^ n16805 ;
  assign n17679 = n16768 ^ n16747 ;
  assign n17678 = n17571 ^ n16768 ;
  assign n17680 = n17679 ^ n17678 ;
  assign n17681 = n17570 & n17680 ;
  assign n17682 = n17681 ^ n17679 ;
  assign n17684 = n17683 ^ n17682 ;
  assign n17685 = n17684 ^ n16768 ;
  assign n17686 = n16039 & ~n17685 ;
  assign n17687 = n17686 ^ n16768 ;
  assign n17673 = n17575 ^ n17564 ;
  assign n17674 = n17575 ^ n15358 ;
  assign n17675 = n17673 & ~n17674 ;
  assign n17676 = n17675 ^ n15358 ;
  assign n17677 = n17676 ^ n15372 ;
  assign n17688 = n17687 ^ n17677 ;
  assign n17690 = n17688 ^ x122 ;
  assign n17689 = n17688 ^ n17576 ;
  assign n17691 = n17690 ^ n17689 ;
  assign n17692 = n17581 & ~n17691 ;
  assign n17693 = n17692 ^ n17690 ;
  assign n17694 = n17693 ^ x121 ;
  assign n17582 = n17581 ^ x122 ;
  assign n17490 = n17489 ^ x123 ;
  assign n17351 = n17350 ^ x124 ;
  assign n17352 = n17268 ^ x113 ;
  assign n17353 = n17262 ^ x114 ;
  assign n17357 = ~n17354 & n17356 ;
  assign n17358 = n17158 ^ x101 ;
  assign n17359 = n17357 & n17358 ;
  assign n17360 = n17165 ^ x100 ;
  assign n17361 = ~n17359 & n17360 ;
  assign n17362 = n17171 ^ x99 ;
  assign n17363 = n17361 & ~n17362 ;
  assign n17364 = n17177 ^ x98 ;
  assign n17365 = n17363 & n17364 ;
  assign n17366 = n17183 ^ x97 ;
  assign n17367 = n17365 & n17366 ;
  assign n17368 = n17189 ^ x96 ;
  assign n17369 = ~n17367 & ~n17368 ;
  assign n17370 = n17195 ^ x111 ;
  assign n17371 = n17369 & n17370 ;
  assign n17372 = n17201 ^ x110 ;
  assign n17373 = ~n17371 & n17372 ;
  assign n17374 = n17206 ^ x109 ;
  assign n17375 = ~n17373 & n17374 ;
  assign n17376 = n17209 ^ x108 ;
  assign n17377 = n17375 & ~n17376 ;
  assign n17378 = n17216 ^ x107 ;
  assign n17379 = ~n17377 & n17378 ;
  assign n17380 = n17223 ^ x106 ;
  assign n17381 = n17379 & n17380 ;
  assign n17382 = n17228 ^ x105 ;
  assign n17383 = n17381 & n17382 ;
  assign n17384 = n17230 ^ n17140 ;
  assign n17385 = n17383 & n17384 ;
  assign n17386 = n17233 ^ x119 ;
  assign n17387 = n17386 ^ n17234 ;
  assign n17388 = ~n17385 & n17387 ;
  assign n17389 = n17240 ^ x118 ;
  assign n17390 = ~n17388 & n17389 ;
  assign n17391 = n17242 ^ x117 ;
  assign n17392 = n17391 ^ n17243 ;
  assign n17393 = ~n17390 & ~n17392 ;
  assign n17394 = n17250 ^ x116 ;
  assign n17395 = ~n17393 & ~n17394 ;
  assign n17396 = n17256 ^ x115 ;
  assign n17397 = ~n17395 & n17396 ;
  assign n17398 = n17353 & ~n17397 ;
  assign n17399 = ~n17352 & ~n17398 ;
  assign n17400 = n17273 ^ x112 ;
  assign n17401 = n17399 & ~n17400 ;
  assign n17402 = n17275 ^ x127 ;
  assign n17403 = n17402 ^ n17290 ;
  assign n17404 = ~n17401 & n17403 ;
  assign n17405 = n17309 ^ x126 ;
  assign n17406 = n17404 & n17405 ;
  assign n17407 = n17329 ^ x125 ;
  assign n17408 = ~n17406 & n17407 ;
  assign n17491 = ~n17351 & ~n17408 ;
  assign n17583 = n17490 & ~n17491 ;
  assign n17672 = n17582 & n17583 ;
  assign n17695 = n17694 ^ n17672 ;
  assign n17584 = n17583 ^ n17582 ;
  assign n17492 = n17491 ^ n17490 ;
  assign n17409 = n17408 ^ n17351 ;
  assign n17410 = n17409 ^ n17015 ;
  assign n17412 = n16891 ^ n16843 ;
  assign n17411 = n17407 ^ n17406 ;
  assign n17413 = n17412 ^ n17411 ;
  assign n17415 = n16886 ^ n16278 ;
  assign n17416 = n17415 ^ n16845 ;
  assign n17414 = n17405 ^ n17404 ;
  assign n17417 = n17416 ^ n17414 ;
  assign n17419 = n16883 ^ n16848 ;
  assign n17420 = n17419 ^ n16847 ;
  assign n17418 = n17403 ^ n17401 ;
  assign n17421 = n17420 ^ n17418 ;
  assign n17423 = n16880 ^ n16246 ;
  assign n17424 = n17423 ^ n16850 ;
  assign n17422 = n17400 ^ n17399 ;
  assign n17425 = n17424 ^ n17422 ;
  assign n17427 = n16878 ^ n16854 ;
  assign n17426 = n17398 ^ n17352 ;
  assign n17428 = n17427 ^ n17426 ;
  assign n17430 = n16874 ^ n16858 ;
  assign n17431 = n17430 ^ n16856 ;
  assign n17429 = n17397 ^ n17353 ;
  assign n17432 = n17431 ^ n17429 ;
  assign n17434 = n16872 ^ n16861 ;
  assign n17433 = n17396 ^ n17395 ;
  assign n17435 = n17434 ^ n17433 ;
  assign n17439 = n16868 ^ n16867 ;
  assign n17436 = n16864 ^ n16863 ;
  assign n17437 = n17392 ^ n17390 ;
  assign n17438 = n17436 & ~n17437 ;
  assign n17440 = n17439 ^ n17438 ;
  assign n17441 = n17394 ^ n17393 ;
  assign n17442 = n17441 ^ n17438 ;
  assign n17443 = ~n17440 & ~n17442 ;
  assign n17444 = n17443 ^ n17439 ;
  assign n17445 = n17444 ^ n17433 ;
  assign n17446 = n17435 & n17445 ;
  assign n17447 = n17446 ^ n17434 ;
  assign n17448 = n17447 ^ n17429 ;
  assign n17449 = n17432 & n17448 ;
  assign n17450 = n17449 ^ n17431 ;
  assign n17451 = n17450 ^ n17426 ;
  assign n17452 = ~n17428 & ~n17451 ;
  assign n17453 = n17452 ^ n17427 ;
  assign n17454 = n17453 ^ n17422 ;
  assign n17455 = ~n17425 & ~n17454 ;
  assign n17456 = n17455 ^ n17424 ;
  assign n17457 = n17456 ^ n17418 ;
  assign n17458 = n17421 & ~n17457 ;
  assign n17459 = n17458 ^ n17420 ;
  assign n17460 = n17459 ^ n17414 ;
  assign n17461 = n17417 & n17460 ;
  assign n17462 = n17461 ^ n17416 ;
  assign n17463 = n17462 ^ n17411 ;
  assign n17464 = n17413 & ~n17463 ;
  assign n17465 = n17464 ^ n17412 ;
  assign n17466 = n17465 ^ n17409 ;
  assign n17467 = ~n17410 & ~n17466 ;
  assign n17468 = n17467 ^ n17015 ;
  assign n17493 = n17492 ^ n17468 ;
  assign n17558 = n17492 ^ n17022 ;
  assign n17559 = n17493 & ~n17558 ;
  assign n17560 = n17559 ^ n17022 ;
  assign n17585 = n17584 ^ n17560 ;
  assign n17669 = n17584 ^ n16954 ;
  assign n17670 = ~n17585 & n17669 ;
  assign n17671 = n17670 ^ n16954 ;
  assign n17696 = n17695 ^ n17671 ;
  assign n17751 = n17695 ^ n16949 ;
  assign n17752 = ~n17696 & ~n17751 ;
  assign n17753 = n17752 ^ n16949 ;
  assign n17744 = n17683 ^ n16768 ;
  assign n17745 = n17682 & n17744 ;
  assign n17742 = n16808 ^ n16807 ;
  assign n17741 = n17683 ^ n16839 ;
  assign n17743 = n17742 ^ n17741 ;
  assign n17746 = n17745 ^ n17743 ;
  assign n17747 = n17746 ^ n16839 ;
  assign n17748 = n16127 & ~n17747 ;
  assign n17738 = n16839 ^ n15388 ;
  assign n17737 = n15372 ^ x120 ;
  assign n17739 = n17738 ^ n17737 ;
  assign n17734 = n17687 ^ n17676 ;
  assign n17735 = n17687 ^ n15372 ;
  assign n17736 = ~n17734 & ~n17735 ;
  assign n17740 = n17739 ^ n17736 ;
  assign n17749 = n17748 ^ n17740 ;
  assign n17729 = n17688 ^ n17672 ;
  assign n17732 = n17693 & ~n17729 ;
  assign n17728 = n17693 ^ n17688 ;
  assign n17730 = n17729 ^ n17728 ;
  assign n17731 = x121 & ~n17730 ;
  assign n17733 = n17732 ^ n17731 ;
  assign n17750 = n17749 ^ n17733 ;
  assign n17754 = n17753 ^ n17750 ;
  assign n17755 = n17753 ^ n16944 ;
  assign n17756 = n17754 & ~n17755 ;
  assign n17757 = n17756 ^ n16944 ;
  assign n17758 = n17757 ^ n17354 ;
  assign n17759 = n17354 ^ n16939 ;
  assign n17760 = ~n17758 & n17759 ;
  assign n17762 = n17761 ^ n17760 ;
  assign n17879 = n17763 ^ n17762 ;
  assign n17873 = n16395 & n17758 ;
  assign n17874 = n17873 ^ n16939 ;
  assign n17863 = n16398 & ~n17754 ;
  assign n17864 = n17863 ^ n16944 ;
  assign n17865 = n17864 ^ n16351 ;
  assign n17697 = ~n16400 & n17696 ;
  assign n17698 = n17697 ^ n16949 ;
  assign n17866 = n17698 ^ n16343 ;
  assign n17586 = ~n16402 & n17585 ;
  assign n17587 = n17586 ^ n16954 ;
  assign n17664 = n17587 ^ n16336 ;
  assign n17494 = ~n16196 & ~n17493 ;
  assign n17495 = n17494 ^ n17022 ;
  assign n17496 = n17495 ^ n16189 ;
  assign n17548 = n16307 & n17466 ;
  assign n17549 = n17548 ^ n17015 ;
  assign n17497 = n16288 & n17463 ;
  assign n17498 = n17497 ^ n17412 ;
  assign n17499 = n17498 ^ n16174 ;
  assign n17500 = n16278 & ~n17460 ;
  assign n17501 = n17500 ^ n17416 ;
  assign n17502 = n17501 ^ n16167 ;
  assign n17503 = n16848 & n17457 ;
  assign n17504 = n17503 ^ n17420 ;
  assign n17505 = n17504 ^ n16164 ;
  assign n17506 = n16246 & n17454 ;
  assign n17507 = n17506 ^ n17424 ;
  assign n17508 = n17507 ^ n15191 ;
  assign n17509 = ~n16853 & n17451 ;
  assign n17510 = n17509 ^ n17427 ;
  assign n17511 = n17510 ^ n16132 ;
  assign n17512 = ~n16858 & ~n17448 ;
  assign n17513 = n17512 ^ n17431 ;
  assign n17514 = n17513 ^ n16137 ;
  assign n17515 = ~n16863 & n17437 ;
  assign n17516 = n17515 ^ n16864 ;
  assign n17517 = ~n16142 & ~n17516 ;
  assign n17518 = n17517 ^ n16145 ;
  assign n17519 = n16866 & n17442 ;
  assign n17520 = n17519 ^ n17439 ;
  assign n17521 = n17520 ^ n17517 ;
  assign n17522 = ~n17518 & n17521 ;
  assign n17523 = n17522 ^ n16145 ;
  assign n17524 = n17523 ^ n16139 ;
  assign n17525 = ~n16860 & ~n17445 ;
  assign n17526 = n17525 ^ n17434 ;
  assign n17527 = n17526 ^ n17523 ;
  assign n17528 = n17524 & n17527 ;
  assign n17529 = n17528 ^ n16139 ;
  assign n17530 = n17529 ^ n17513 ;
  assign n17531 = ~n17514 & ~n17530 ;
  assign n17532 = n17531 ^ n16137 ;
  assign n17533 = n17532 ^ n17510 ;
  assign n17534 = n17511 & ~n17533 ;
  assign n17535 = n17534 ^ n16132 ;
  assign n17536 = n17535 ^ n17507 ;
  assign n17537 = ~n17508 & n17536 ;
  assign n17538 = n17537 ^ n15191 ;
  assign n17539 = n17538 ^ n17504 ;
  assign n17540 = n17505 & n17539 ;
  assign n17541 = n17540 ^ n16164 ;
  assign n17542 = n17541 ^ n17501 ;
  assign n17543 = n17502 & n17542 ;
  assign n17544 = n17543 ^ n16167 ;
  assign n17545 = n17544 ^ n17498 ;
  assign n17546 = n17499 & ~n17545 ;
  assign n17547 = n17546 ^ n16174 ;
  assign n17550 = n17549 ^ n17547 ;
  assign n17551 = n17549 ^ n16182 ;
  assign n17552 = n17550 & n17551 ;
  assign n17553 = n17552 ^ n16182 ;
  assign n17554 = n17553 ^ n17495 ;
  assign n17555 = ~n17496 & ~n17554 ;
  assign n17556 = n17555 ^ n16189 ;
  assign n17665 = n17587 ^ n17556 ;
  assign n17666 = ~n17664 & n17665 ;
  assign n17667 = n17666 ^ n16336 ;
  assign n17867 = n17698 ^ n17667 ;
  assign n17868 = n17866 & ~n17867 ;
  assign n17869 = n17868 ^ n16343 ;
  assign n17870 = n17869 ^ n17864 ;
  assign n17871 = n17865 & n17870 ;
  assign n17872 = n17871 ^ n16351 ;
  assign n17875 = n17874 ^ n17872 ;
  assign n17876 = n17874 ^ n16358 ;
  assign n17877 = ~n17875 & n17876 ;
  assign n17878 = n17877 ^ n16358 ;
  assign n18035 = n17878 ^ n16366 ;
  assign n17880 = n17879 ^ n17042 ;
  assign n17881 = n16396 & ~n17880 ;
  assign n17882 = n17881 ^ n17042 ;
  assign n18036 = n18035 ^ n17882 ;
  assign n18016 = n17872 ^ n16358 ;
  assign n18017 = n18016 ^ n17874 ;
  assign n18018 = n18017 ^ x265 ;
  assign n17668 = n17667 ^ n16343 ;
  assign n17699 = n17698 ^ n17668 ;
  assign n17557 = n17556 ^ n16336 ;
  assign n17588 = n17587 ^ n17557 ;
  assign n17589 = n17588 ^ x268 ;
  assign n17591 = n17516 ^ n16142 ;
  assign n17592 = x263 & n17591 ;
  assign n17590 = n17520 ^ n17518 ;
  assign n17593 = n17592 ^ n17590 ;
  assign n17594 = n17526 ^ n17524 ;
  assign n17595 = n17594 ^ x262 ;
  assign n17596 = n17595 ^ n17590 ;
  assign n17597 = n17596 ^ n17594 ;
  assign n17598 = ~n17593 & n17597 ;
  assign n17599 = n17598 ^ n17595 ;
  assign n17600 = n17529 ^ n16137 ;
  assign n17601 = n17600 ^ n17513 ;
  assign n17603 = n17601 ^ x261 ;
  assign n17602 = n17601 ^ n17594 ;
  assign n17604 = n17603 ^ n17602 ;
  assign n17605 = ~n17599 & n17604 ;
  assign n17606 = n17605 ^ n17603 ;
  assign n17607 = n17532 ^ n16132 ;
  assign n17608 = n17607 ^ n17510 ;
  assign n17610 = n17608 ^ x260 ;
  assign n17609 = n17608 ^ n17601 ;
  assign n17611 = n17610 ^ n17609 ;
  assign n17612 = ~n17606 & n17611 ;
  assign n17613 = n17612 ^ n17610 ;
  assign n17614 = n17535 ^ n15191 ;
  assign n17615 = n17614 ^ n17507 ;
  assign n17617 = n17615 ^ x259 ;
  assign n17616 = n17615 ^ n17608 ;
  assign n17618 = n17617 ^ n17616 ;
  assign n17619 = ~n17613 & n17618 ;
  assign n17620 = n17619 ^ n17617 ;
  assign n17621 = n17538 ^ n16164 ;
  assign n17622 = n17621 ^ n17504 ;
  assign n17624 = n17622 ^ x258 ;
  assign n17623 = n17622 ^ n17615 ;
  assign n17625 = n17624 ^ n17623 ;
  assign n17626 = n17620 & ~n17625 ;
  assign n17627 = n17626 ^ n17624 ;
  assign n17628 = n17541 ^ n16167 ;
  assign n17629 = n17628 ^ n17501 ;
  assign n17631 = n17629 ^ x257 ;
  assign n17630 = n17629 ^ n17622 ;
  assign n17632 = n17631 ^ n17630 ;
  assign n17633 = ~n17627 & n17632 ;
  assign n17634 = n17633 ^ n17631 ;
  assign n17635 = n17544 ^ n16174 ;
  assign n17636 = n17635 ^ n17498 ;
  assign n17638 = n17636 ^ x256 ;
  assign n17637 = n17636 ^ n17629 ;
  assign n17639 = n17638 ^ n17637 ;
  assign n17640 = n17634 & ~n17639 ;
  assign n17641 = n17640 ^ n17638 ;
  assign n17642 = n17547 ^ n16182 ;
  assign n17643 = n17642 ^ n17549 ;
  assign n17645 = n17643 ^ x271 ;
  assign n17644 = n17643 ^ n17636 ;
  assign n17646 = n17645 ^ n17644 ;
  assign n17647 = ~n17641 & n17646 ;
  assign n17648 = n17647 ^ n17645 ;
  assign n17649 = n17553 ^ n16189 ;
  assign n17650 = n17649 ^ n17495 ;
  assign n17652 = n17650 ^ x270 ;
  assign n17651 = n17650 ^ n17643 ;
  assign n17653 = n17652 ^ n17651 ;
  assign n17654 = ~n17648 & n17653 ;
  assign n17655 = n17654 ^ n17652 ;
  assign n17657 = n17588 ^ x269 ;
  assign n17656 = n17650 ^ n17588 ;
  assign n17658 = n17657 ^ n17656 ;
  assign n17659 = ~n17655 & n17658 ;
  assign n17660 = n17659 ^ n17657 ;
  assign n17661 = ~n17589 & n17660 ;
  assign n17662 = n17661 ^ x268 ;
  assign n18019 = n17699 ^ n17662 ;
  assign n18020 = n17869 ^ n16351 ;
  assign n18021 = n18020 ^ n17864 ;
  assign n18022 = n18021 ^ x267 ;
  assign n18023 = n18022 ^ n17662 ;
  assign n18024 = n18023 ^ n18021 ;
  assign n18025 = ~n18019 & n18024 ;
  assign n18026 = n18025 ^ n18022 ;
  assign n18028 = n18017 ^ x266 ;
  assign n18027 = n18021 ^ n18017 ;
  assign n18029 = n18028 ^ n18027 ;
  assign n18030 = ~n18026 & n18029 ;
  assign n18031 = n18030 ^ n18028 ;
  assign n18032 = ~n18018 & n18031 ;
  assign n18033 = n18032 ^ x265 ;
  assign n18037 = n18036 ^ n18033 ;
  assign n18146 = n18037 ^ x264 ;
  assign n17663 = n17662 ^ x267 ;
  assign n17700 = n17699 ^ n17663 ;
  assign n17701 = n17591 ^ x263 ;
  assign n17702 = n17592 ^ x262 ;
  assign n17703 = n17702 ^ n17590 ;
  assign n17704 = n17701 & n17703 ;
  assign n17705 = n17599 ^ x261 ;
  assign n17706 = ~n17704 & ~n17705 ;
  assign n17707 = n17606 ^ x260 ;
  assign n17708 = n17706 & ~n17707 ;
  assign n17709 = n17613 ^ x259 ;
  assign n17710 = ~n17708 & n17709 ;
  assign n17711 = n17620 ^ x258 ;
  assign n17712 = ~n17710 & n17711 ;
  assign n17713 = n17627 ^ x257 ;
  assign n17714 = n17712 & ~n17713 ;
  assign n17715 = n17634 ^ x256 ;
  assign n17716 = n17714 & n17715 ;
  assign n17717 = n17641 ^ x271 ;
  assign n17718 = ~n17716 & n17717 ;
  assign n17719 = n17648 ^ x270 ;
  assign n17720 = n17718 & n17719 ;
  assign n17721 = n17655 ^ x269 ;
  assign n17722 = ~n17720 & ~n17721 ;
  assign n17723 = n17660 ^ x268 ;
  assign n17724 = ~n17722 & ~n17723 ;
  assign n18141 = ~n17700 & ~n17724 ;
  assign n18142 = n18026 ^ x266 ;
  assign n18143 = ~n18141 & n18142 ;
  assign n18144 = n18031 ^ x265 ;
  assign n18145 = n18143 & ~n18144 ;
  assign n18213 = n18146 ^ n18145 ;
  assign n18211 = n17447 ^ n17431 ;
  assign n18212 = n18211 ^ n17429 ;
  assign n18214 = n18213 ^ n18212 ;
  assign n18216 = n17444 ^ n17434 ;
  assign n18217 = n18216 ^ n17433 ;
  assign n18215 = n18144 ^ n18143 ;
  assign n18218 = n18217 ^ n18215 ;
  assign n18220 = n17441 ^ n17440 ;
  assign n17725 = n17724 ^ n17700 ;
  assign n17726 = n17437 ^ n17436 ;
  assign n18219 = ~n17725 & ~n17726 ;
  assign n18221 = n18220 ^ n18219 ;
  assign n18222 = n18142 ^ n18141 ;
  assign n18223 = n18222 ^ n18219 ;
  assign n18224 = ~n18221 & n18223 ;
  assign n18225 = n18224 ^ n18220 ;
  assign n18226 = n18225 ^ n18215 ;
  assign n18227 = n18218 & ~n18226 ;
  assign n18228 = n18227 ^ n18217 ;
  assign n18229 = n18228 ^ n18212 ;
  assign n18230 = ~n18214 & n18229 ;
  assign n18231 = n18230 ^ n18213 ;
  assign n18147 = n18145 & ~n18146 ;
  assign n18034 = n18033 ^ x264 ;
  assign n18038 = n18034 & n18037 ;
  assign n18039 = n18038 ^ x264 ;
  assign n18139 = n18039 ^ x279 ;
  assign n17883 = n17882 ^ n17878 ;
  assign n17770 = n17358 ^ n17357 ;
  assign n17765 = n17047 ^ n17042 ;
  assign n17764 = n17763 ^ n17047 ;
  assign n17766 = n17765 ^ n17764 ;
  assign n17767 = n17762 & ~n17766 ;
  assign n17768 = n17767 ^ n17765 ;
  assign n17858 = n17770 ^ n17768 ;
  assign n17859 = n17858 ^ n17047 ;
  assign n17860 = n16919 & n17859 ;
  assign n17861 = n17860 ^ n17047 ;
  assign n17884 = n17861 ^ n16366 ;
  assign n17885 = n17884 ^ n17861 ;
  assign n17886 = n17885 ^ n17878 ;
  assign n17887 = ~n17883 & n17886 ;
  assign n17888 = n17887 ^ n17884 ;
  assign n18015 = n17888 ^ n16378 ;
  assign n18140 = n18139 ^ n18015 ;
  assign n18207 = n18147 ^ n18140 ;
  assign n18232 = n18231 ^ n18207 ;
  assign n18312 = n17427 & n18232 ;
  assign n18208 = n17450 ^ n17427 ;
  assign n18209 = n18208 ^ n17426 ;
  assign n18313 = n18312 ^ n18209 ;
  assign n18314 = n18313 ^ n16853 ;
  assign n18315 = n17434 & n18226 ;
  assign n18316 = n18315 ^ n18217 ;
  assign n18317 = n18316 ^ n16860 ;
  assign n18318 = n17436 & n17725 ;
  assign n18319 = n18318 ^ n17437 ;
  assign n18320 = ~n16863 & ~n18319 ;
  assign n18321 = n18320 ^ n16866 ;
  assign n18322 = ~n17439 & ~n18223 ;
  assign n18323 = n18322 ^ n18220 ;
  assign n18324 = n18323 ^ n18320 ;
  assign n18325 = n18321 & n18324 ;
  assign n18326 = n18325 ^ n16866 ;
  assign n18327 = n18326 ^ n18316 ;
  assign n18328 = n18317 & n18327 ;
  assign n18329 = n18328 ^ n16860 ;
  assign n18330 = n18329 ^ n16858 ;
  assign n18331 = n18228 ^ n18213 ;
  assign n18332 = ~n17431 & n18331 ;
  assign n18333 = n18332 ^ n18212 ;
  assign n18334 = n18333 ^ n18329 ;
  assign n18335 = n18330 & n18334 ;
  assign n18336 = n18335 ^ n16858 ;
  assign n18337 = n18336 ^ n18313 ;
  assign n18338 = ~n18314 & n18337 ;
  assign n18339 = n18338 ^ n16853 ;
  assign n18495 = n18339 ^ n16246 ;
  assign n18210 = n18209 ^ n18207 ;
  assign n18233 = ~n18210 & ~n18232 ;
  assign n18234 = n18233 ^ n18209 ;
  assign n18148 = ~n18140 & n18147 ;
  assign n18040 = n18039 ^ n18015 ;
  assign n17862 = n17861 ^ n16378 ;
  assign n17889 = n17862 & n17888 ;
  assign n17890 = n17889 ^ n16378 ;
  assign n18041 = n17890 ^ n16384 ;
  assign n17769 = n17360 ^ n17359 ;
  assign n17772 = n17769 ^ n17047 ;
  assign n17771 = n17770 ^ n17769 ;
  assign n17773 = n17772 ^ n17771 ;
  assign n17774 = ~n17768 & ~n17773 ;
  assign n17775 = n17774 ^ n17772 ;
  assign n17891 = ~n16385 & ~n17775 ;
  assign n17892 = n17891 ^ n17059 ;
  assign n18042 = n18041 ^ n17892 ;
  assign n18043 = n18042 ^ x279 ;
  assign n18044 = n18043 ^ n18015 ;
  assign n18045 = n18044 ^ n18042 ;
  assign n18046 = n18040 & ~n18045 ;
  assign n18047 = n18046 ^ n18043 ;
  assign n18138 = n18047 ^ x278 ;
  assign n18205 = n18148 ^ n18138 ;
  assign n18340 = n18234 ^ n18205 ;
  assign n18341 = ~n17424 & n18340 ;
  assign n18203 = n17453 ^ n17424 ;
  assign n18204 = n18203 ^ n17422 ;
  assign n18342 = n18341 ^ n18204 ;
  assign n18496 = n18495 ^ n18342 ;
  assign n18497 = n18496 ^ x418 ;
  assign n18513 = n18333 ^ n18330 ;
  assign n18500 = n18319 ^ n16863 ;
  assign n18501 = x423 & n18500 ;
  assign n18502 = n18501 ^ x422 ;
  assign n18503 = n18323 ^ n18321 ;
  assign n18504 = n18503 ^ n18501 ;
  assign n18505 = n18502 & n18504 ;
  assign n18506 = n18505 ^ x422 ;
  assign n18507 = n18506 ^ x421 ;
  assign n18508 = n18326 ^ n16860 ;
  assign n18509 = n18508 ^ n18316 ;
  assign n18510 = n18509 ^ n18506 ;
  assign n18511 = n18507 & ~n18510 ;
  assign n18512 = n18511 ^ x421 ;
  assign n18514 = n18513 ^ n18512 ;
  assign n18515 = n18512 ^ x420 ;
  assign n18516 = ~n18514 & n18515 ;
  assign n18517 = n18516 ^ x420 ;
  assign n18498 = n18336 ^ n16853 ;
  assign n18499 = n18498 ^ n18313 ;
  assign n18518 = n18517 ^ n18499 ;
  assign n18520 = n18496 ^ x419 ;
  assign n18519 = n18517 ^ n18496 ;
  assign n18521 = n18520 ^ n18519 ;
  assign n18522 = ~n18518 & n18521 ;
  assign n18523 = n18522 ^ n18520 ;
  assign n18524 = n18497 & ~n18523 ;
  assign n18525 = n18524 ^ x418 ;
  assign n18343 = n18342 ^ n18339 ;
  assign n18344 = n18342 ^ n16246 ;
  assign n18345 = ~n18343 & ~n18344 ;
  assign n18346 = n18345 ^ n16246 ;
  assign n18493 = n18346 ^ n16848 ;
  assign n18206 = n18205 ^ n18204 ;
  assign n18235 = n18234 ^ n18204 ;
  assign n18236 = ~n18206 & n18235 ;
  assign n18237 = n18236 ^ n18205 ;
  assign n18149 = n18138 & ~n18148 ;
  assign n17893 = n17892 ^ n17890 ;
  assign n17894 = n17892 ^ n16384 ;
  assign n17895 = n17893 & ~n17894 ;
  assign n17896 = n17895 ^ n16384 ;
  assign n18048 = n17896 ^ n16198 ;
  assign n17782 = n17362 ^ n17361 ;
  assign n17777 = n17059 ^ n16934 ;
  assign n17776 = n17769 ^ n16934 ;
  assign n17778 = n17777 ^ n17776 ;
  assign n17779 = n17775 & n17778 ;
  assign n17780 = n17779 ^ n17777 ;
  assign n17897 = n17782 ^ n17780 ;
  assign n17898 = n17897 ^ n16934 ;
  assign n17899 = ~n16391 & n17898 ;
  assign n17900 = n17899 ^ n16934 ;
  assign n18049 = n18048 ^ n17900 ;
  assign n18051 = n18049 ^ x278 ;
  assign n18050 = n18049 ^ n18042 ;
  assign n18052 = n18051 ^ n18050 ;
  assign n18053 = n18047 & ~n18052 ;
  assign n18054 = n18053 ^ n18051 ;
  assign n18137 = n18054 ^ x277 ;
  assign n18201 = n18149 ^ n18137 ;
  assign n18347 = n18237 ^ n18201 ;
  assign n18348 = ~n17420 & ~n18347 ;
  assign n18199 = n17456 ^ n17420 ;
  assign n18200 = n18199 ^ n17418 ;
  assign n18349 = n18348 ^ n18200 ;
  assign n18494 = n18493 ^ n18349 ;
  assign n18526 = n18525 ^ n18494 ;
  assign n18527 = n18525 ^ x417 ;
  assign n18528 = n18526 & n18527 ;
  assign n18529 = n18528 ^ x417 ;
  assign n18350 = n18349 ^ n18346 ;
  assign n18351 = n18349 ^ n16848 ;
  assign n18352 = n18350 & ~n18351 ;
  assign n18353 = n18352 ^ n16848 ;
  assign n18491 = n18353 ^ n16278 ;
  assign n18202 = n18201 ^ n18200 ;
  assign n18238 = n18237 ^ n18200 ;
  assign n18239 = n18202 & n18238 ;
  assign n18240 = n18239 ^ n18201 ;
  assign n18150 = n18137 & ~n18149 ;
  assign n17901 = n17900 ^ n17896 ;
  assign n17902 = n17900 ^ n16198 ;
  assign n17903 = ~n17901 & n17902 ;
  assign n17904 = n17903 ^ n16198 ;
  assign n18055 = n17904 ^ n16407 ;
  assign n17781 = n17364 ^ n17363 ;
  assign n17784 = n17781 ^ n16934 ;
  assign n17783 = n17782 ^ n17781 ;
  assign n17785 = n17784 ^ n17783 ;
  assign n17786 = ~n17780 & ~n17785 ;
  assign n17787 = n17786 ^ n17784 ;
  assign n17905 = n16444 & n17787 ;
  assign n17906 = n17905 ^ n17077 ;
  assign n18056 = n18055 ^ n17906 ;
  assign n18058 = n18056 ^ x277 ;
  assign n18057 = n18056 ^ n18049 ;
  assign n18059 = n18058 ^ n18057 ;
  assign n18060 = ~n18054 & n18059 ;
  assign n18061 = n18060 ^ n18058 ;
  assign n18136 = n18061 ^ x276 ;
  assign n18197 = n18150 ^ n18136 ;
  assign n18308 = n18240 ^ n18197 ;
  assign n18309 = n17416 & n18308 ;
  assign n18195 = n17459 ^ n17416 ;
  assign n18196 = n18195 ^ n17414 ;
  assign n18310 = n18309 ^ n18196 ;
  assign n18492 = n18491 ^ n18310 ;
  assign n18530 = n18529 ^ n18492 ;
  assign n18198 = n18197 ^ n18196 ;
  assign n18241 = n18240 ^ n18196 ;
  assign n18242 = n18198 & ~n18241 ;
  assign n18243 = n18242 ^ n18197 ;
  assign n18151 = ~n18136 & ~n18150 ;
  assign n17907 = n17906 ^ n17904 ;
  assign n17908 = n17906 ^ n16407 ;
  assign n17909 = ~n17907 & n17908 ;
  assign n17910 = n17909 ^ n16407 ;
  assign n18062 = n17910 ^ n15624 ;
  assign n17798 = n17366 ^ n17365 ;
  assign n17794 = n17090 ^ n17077 ;
  assign n17793 = n17781 ^ n17090 ;
  assign n17795 = n17794 ^ n17793 ;
  assign n17796 = ~n17787 & n17795 ;
  assign n17797 = n17796 ^ n17794 ;
  assign n17911 = n17798 ^ n17797 ;
  assign n17912 = n17911 ^ n17090 ;
  assign n17913 = n16439 & n17912 ;
  assign n17914 = n17913 ^ n17090 ;
  assign n18063 = n18062 ^ n17914 ;
  assign n18065 = n18063 ^ x276 ;
  assign n18064 = n18063 ^ n18056 ;
  assign n18066 = n18065 ^ n18064 ;
  assign n18067 = ~n18061 & n18066 ;
  assign n18068 = n18067 ^ n18065 ;
  assign n18135 = n18068 ^ x275 ;
  assign n18194 = n18151 ^ n18135 ;
  assign n18244 = n18243 ^ n18194 ;
  assign n18358 = n17412 & ~n18244 ;
  assign n18245 = n17462 ^ n17412 ;
  assign n18246 = n18245 ^ n17411 ;
  assign n18359 = n18358 ^ n18246 ;
  assign n18311 = n18310 ^ n16278 ;
  assign n18354 = n18353 ^ n18310 ;
  assign n18355 = ~n18311 & n18354 ;
  assign n18356 = n18355 ^ n16278 ;
  assign n18357 = n18356 ^ n16288 ;
  assign n18531 = n18359 ^ n18357 ;
  assign n18532 = n18531 ^ x416 ;
  assign n18533 = n18532 ^ n18529 ;
  assign n18534 = n18533 ^ n18531 ;
  assign n18535 = n18530 & n18534 ;
  assign n18536 = n18535 ^ n18532 ;
  assign n18247 = n18246 ^ n18194 ;
  assign n18248 = ~n18244 & ~n18247 ;
  assign n18249 = n18248 ^ n18243 ;
  assign n18152 = ~n18135 & n18151 ;
  assign n17915 = n17914 ^ n17910 ;
  assign n17804 = n17368 ^ n17367 ;
  assign n17800 = n17103 ^ n17090 ;
  assign n17799 = n17798 ^ n17103 ;
  assign n17801 = n17800 ^ n17799 ;
  assign n17802 = ~n17797 & ~n17801 ;
  assign n17803 = n17802 ^ n17800 ;
  assign n17853 = n17804 ^ n17803 ;
  assign n17854 = n17853 ^ n17103 ;
  assign n17855 = n16434 & n17854 ;
  assign n17856 = n17855 ^ n17103 ;
  assign n17916 = n17856 ^ n15624 ;
  assign n17917 = n17916 ^ n17856 ;
  assign n17918 = n17917 ^ n17910 ;
  assign n17919 = n17915 & ~n17918 ;
  assign n17920 = n17919 ^ n17916 ;
  assign n18069 = n17920 ^ n15619 ;
  assign n18071 = n18069 ^ x275 ;
  assign n18070 = n18069 ^ n18063 ;
  assign n18072 = n18071 ^ n18070 ;
  assign n18073 = ~n18068 & n18072 ;
  assign n18074 = n18073 ^ n18071 ;
  assign n18134 = n18074 ^ x274 ;
  assign n18192 = n18152 ^ n18134 ;
  assign n18364 = n18249 ^ n18192 ;
  assign n18365 = ~n17015 & ~n18364 ;
  assign n18190 = n17465 ^ n17015 ;
  assign n18191 = n18190 ^ n17409 ;
  assign n18366 = n18365 ^ n18191 ;
  assign n18360 = n18359 ^ n18356 ;
  assign n18361 = n18357 & ~n18360 ;
  assign n18362 = n18361 ^ n16288 ;
  assign n18363 = n18362 ^ n16307 ;
  assign n18537 = n18366 ^ n18363 ;
  assign n18539 = n18537 ^ x431 ;
  assign n18538 = n18537 ^ n18531 ;
  assign n18540 = n18539 ^ n18538 ;
  assign n18541 = ~n18536 & n18540 ;
  assign n18542 = n18541 ^ n18539 ;
  assign n18193 = n18192 ^ n18191 ;
  assign n18250 = n18249 ^ n18191 ;
  assign n18251 = ~n18193 & ~n18250 ;
  assign n18252 = n18251 ^ n18192 ;
  assign n17857 = n17856 ^ n15619 ;
  assign n17921 = n17857 & ~n17920 ;
  assign n17922 = n17921 ^ n15619 ;
  assign n18075 = n17922 ^ n15761 ;
  assign n17810 = n17370 ^ n17369 ;
  assign n17806 = n17116 ^ n17103 ;
  assign n17805 = n17804 ^ n17116 ;
  assign n17807 = n17806 ^ n17805 ;
  assign n17808 = n17803 & n17807 ;
  assign n17809 = n17808 ^ n17806 ;
  assign n17923 = n17810 ^ n17809 ;
  assign n17924 = n17923 ^ n17116 ;
  assign n17925 = n16429 & n17924 ;
  assign n17926 = n17925 ^ n17116 ;
  assign n18076 = n18075 ^ n17926 ;
  assign n18078 = n18076 ^ x274 ;
  assign n18077 = n18076 ^ n18069 ;
  assign n18079 = n18078 ^ n18077 ;
  assign n18080 = n18074 & ~n18079 ;
  assign n18081 = n18080 ^ n18078 ;
  assign n18154 = n18081 ^ x273 ;
  assign n18153 = ~n18134 & ~n18152 ;
  assign n18188 = n18154 ^ n18153 ;
  assign n18371 = n18252 ^ n18188 ;
  assign n18372 = ~n17022 & n18371 ;
  assign n18186 = n17468 ^ n17022 ;
  assign n18187 = n18186 ^ n17492 ;
  assign n18373 = n18372 ^ n18187 ;
  assign n18367 = n18366 ^ n18362 ;
  assign n18368 = n18363 & n18367 ;
  assign n18369 = n18368 ^ n16307 ;
  assign n18370 = n18369 ^ n16196 ;
  assign n18543 = n18373 ^ n18370 ;
  assign n18545 = n18543 ^ x430 ;
  assign n18544 = n18543 ^ n18537 ;
  assign n18546 = n18545 ^ n18544 ;
  assign n18547 = n18542 & ~n18546 ;
  assign n18548 = n18547 ^ n18545 ;
  assign n18704 = n18548 ^ x429 ;
  assign n18684 = n18526 ^ x417 ;
  assign n18685 = n16863 ^ x423 ;
  assign n18686 = n18685 ^ n18319 ;
  assign n18687 = n18504 ^ x422 ;
  assign n18688 = n18686 & ~n18687 ;
  assign n18689 = n18510 ^ x421 ;
  assign n18690 = ~n18688 & ~n18689 ;
  assign n18691 = n18514 ^ x420 ;
  assign n18692 = ~n18690 & n18691 ;
  assign n18693 = n18518 ^ x419 ;
  assign n18694 = n18692 & n18693 ;
  assign n18695 = n18523 ^ x418 ;
  assign n18696 = n18694 & n18695 ;
  assign n18697 = ~n18684 & n18696 ;
  assign n18698 = n18530 ^ x416 ;
  assign n18699 = n18697 & ~n18698 ;
  assign n18700 = n18536 ^ x431 ;
  assign n18701 = ~n18699 & ~n18700 ;
  assign n18702 = n18542 ^ x430 ;
  assign n18703 = ~n18701 & ~n18702 ;
  assign n18973 = n18704 ^ n18703 ;
  assign n17927 = n17926 ^ n17922 ;
  assign n17928 = n17926 ^ n15761 ;
  assign n17929 = ~n17927 & n17928 ;
  assign n17930 = n17929 ^ n15761 ;
  assign n18012 = n17930 ^ n16529 ;
  assign n17816 = n17372 ^ n17371 ;
  assign n17812 = n17129 ^ n17116 ;
  assign n17811 = n17810 ^ n17129 ;
  assign n17813 = n17812 ^ n17811 ;
  assign n17814 = n17809 & n17813 ;
  assign n17815 = n17814 ^ n17812 ;
  assign n17931 = n17816 ^ n17815 ;
  assign n17932 = n17931 ^ n17129 ;
  assign n17933 = n16536 & n17932 ;
  assign n17934 = n17933 ^ n17129 ;
  assign n18013 = n18012 ^ n17934 ;
  assign n18014 = n18013 ^ x272 ;
  assign n18083 = n18013 ^ x273 ;
  assign n18082 = n18076 ^ n18013 ;
  assign n18084 = n18083 ^ n18082 ;
  assign n18085 = n18081 & ~n18084 ;
  assign n18086 = n18085 ^ n18083 ;
  assign n18087 = n18014 & ~n18086 ;
  assign n18088 = n18087 ^ x272 ;
  assign n17935 = n17934 ^ n17930 ;
  assign n17791 = n17282 ^ n16645 ;
  assign n17818 = n17791 ^ n17129 ;
  assign n17817 = n17816 ^ n17791 ;
  assign n17819 = n17818 ^ n17817 ;
  assign n17820 = n17815 & n17819 ;
  assign n17821 = n17820 ^ n17818 ;
  assign n17790 = n17374 ^ n17373 ;
  assign n17848 = n17821 ^ n17790 ;
  assign n17849 = n17848 ^ n17282 ;
  assign n17850 = n16645 & n17849 ;
  assign n17851 = n17850 ^ n17848 ;
  assign n17936 = n17851 ^ n16529 ;
  assign n17937 = n17936 ^ n17930 ;
  assign n17938 = n17937 ^ n17851 ;
  assign n17939 = ~n17935 & ~n17938 ;
  assign n17940 = n17939 ^ n17936 ;
  assign n18011 = n17940 ^ n16638 ;
  assign n18089 = n18088 ^ n18011 ;
  assign n17792 = n17791 ^ n17790 ;
  assign n17822 = ~n17792 & n17821 ;
  assign n17823 = n17822 ^ n17791 ;
  assign n17789 = n17376 ^ n17375 ;
  assign n17824 = n17823 ^ n17789 ;
  assign n17944 = ~n17314 & n17824 ;
  assign n17945 = n17944 ^ n17296 ;
  assign n17852 = n17851 ^ n16638 ;
  assign n17941 = ~n17852 & ~n17940 ;
  assign n17942 = n17941 ^ n16638 ;
  assign n17943 = n17942 ^ n16678 ;
  assign n18090 = n17945 ^ n17943 ;
  assign n18091 = n18090 ^ x287 ;
  assign n18092 = n18091 ^ n18011 ;
  assign n18093 = n18092 ^ n18090 ;
  assign n18094 = n18089 & ~n18093 ;
  assign n18095 = n18094 ^ n18091 ;
  assign n18131 = n18095 ^ x286 ;
  assign n18132 = n18088 ^ x287 ;
  assign n18133 = n18132 ^ n18011 ;
  assign n18155 = ~n18153 & n18154 ;
  assign n18156 = n18086 ^ x272 ;
  assign n18157 = ~n18155 & n18156 ;
  assign n18158 = n18133 & ~n18157 ;
  assign n18159 = n18131 & ~n18158 ;
  assign n17946 = n17945 ^ n17942 ;
  assign n17947 = n17943 & n17946 ;
  assign n17948 = n17947 ^ n16678 ;
  assign n18008 = n17948 ^ n15952 ;
  assign n17830 = n17378 ^ n17377 ;
  assign n17828 = n17789 ^ n17320 ;
  assign n17825 = n17314 ^ n17296 ;
  assign n17826 = n17825 ^ n17789 ;
  assign n17827 = ~n17824 & ~n17826 ;
  assign n17829 = n17828 ^ n17827 ;
  assign n17949 = n17830 ^ n17829 ;
  assign n17950 = n17949 ^ n17320 ;
  assign n17951 = ~n16684 & ~n17950 ;
  assign n17952 = n17951 ^ n17320 ;
  assign n18009 = n18008 ^ n17952 ;
  assign n18097 = n18009 ^ x286 ;
  assign n18096 = n18090 ^ n18009 ;
  assign n18098 = n18097 ^ n18096 ;
  assign n18099 = ~n18095 & n18098 ;
  assign n18100 = n18099 ^ n18097 ;
  assign n18130 = n18100 ^ x285 ;
  assign n18178 = n18159 ^ n18130 ;
  assign n18177 = n17759 ^ n17757 ;
  assign n18179 = n18178 ^ n18177 ;
  assign n18183 = n18157 ^ n18133 ;
  assign n18181 = n17671 ^ n16949 ;
  assign n18182 = n18181 ^ n17695 ;
  assign n18184 = n18183 ^ n18182 ;
  assign n18189 = n18188 ^ n18187 ;
  assign n18253 = n18252 ^ n18187 ;
  assign n18254 = n18189 & ~n18253 ;
  assign n18255 = n18254 ^ n18188 ;
  assign n18185 = n18156 ^ n18155 ;
  assign n18256 = n18255 ^ n18185 ;
  assign n18257 = n17560 ^ n16954 ;
  assign n18258 = n18257 ^ n17584 ;
  assign n18259 = n18258 ^ n18185 ;
  assign n18260 = ~n18256 & ~n18259 ;
  assign n18261 = n18260 ^ n18255 ;
  assign n18262 = n18261 ^ n18182 ;
  assign n18263 = n18184 & ~n18262 ;
  assign n18264 = n18263 ^ n18183 ;
  assign n18180 = n18158 ^ n18131 ;
  assign n18265 = n18264 ^ n18180 ;
  assign n18266 = n17755 ^ n17750 ;
  assign n18267 = n18266 ^ n18180 ;
  assign n18268 = ~n18265 & n18267 ;
  assign n18269 = n18268 ^ n18264 ;
  assign n18270 = n18269 ^ n18177 ;
  assign n18271 = ~n18179 & n18270 ;
  assign n18272 = n18271 ^ n18178 ;
  assign n18969 = n18272 ^ n17879 ;
  assign n18160 = n18130 & ~n18159 ;
  assign n17953 = n17952 ^ n17948 ;
  assign n17954 = n17952 ^ n15952 ;
  assign n17955 = n17953 & n17954 ;
  assign n17956 = n17955 ^ n15952 ;
  assign n18103 = n17956 ^ n15976 ;
  assign n17836 = n17380 ^ n17379 ;
  assign n17832 = n17341 ^ n17320 ;
  assign n17831 = n17830 ^ n17341 ;
  assign n17833 = n17832 ^ n17831 ;
  assign n17834 = n17829 & ~n17833 ;
  assign n17835 = n17834 ^ n17832 ;
  assign n17957 = n17836 ^ n17835 ;
  assign n17958 = n17957 ^ n17341 ;
  assign n17959 = n16705 & n17958 ;
  assign n17960 = n17959 ^ n17341 ;
  assign n18104 = n18103 ^ n17960 ;
  assign n18128 = n18104 ^ x284 ;
  assign n18010 = n18009 ^ x285 ;
  assign n18101 = ~n18010 & n18100 ;
  assign n18102 = n18101 ^ x285 ;
  assign n18129 = n18128 ^ n18102 ;
  assign n18273 = n18160 ^ n18129 ;
  assign n18970 = n18969 ^ n18273 ;
  assign n18770 = n18270 ^ n18178 ;
  assign n18971 = n18970 ^ n18770 ;
  assign n18774 = n18250 ^ n18192 ;
  assign n18771 = n18693 ^ n18692 ;
  assign n18775 = n18774 ^ n18771 ;
  assign n18779 = n18691 ^ n18690 ;
  assign n18776 = n18246 ^ n18243 ;
  assign n18777 = n18776 ^ n18194 ;
  assign n18780 = n18779 ^ n18777 ;
  assign n18868 = n18235 ^ n18205 ;
  assign n18646 = n17825 ^ n17824 ;
  assign n18105 = n18104 ^ n18102 ;
  assign n17961 = n17960 ^ n17956 ;
  assign n17962 = n17960 ^ n15976 ;
  assign n17963 = ~n17961 & n17962 ;
  assign n17964 = n17963 ^ n15976 ;
  assign n17842 = n17382 ^ n17381 ;
  assign n17838 = n17480 ^ n17341 ;
  assign n17837 = n17836 ^ n17480 ;
  assign n17839 = n17838 ^ n17837 ;
  assign n17840 = n17835 & n17839 ;
  assign n17841 = n17840 ^ n17838 ;
  assign n17843 = n17842 ^ n17841 ;
  assign n17844 = n17843 ^ n17480 ;
  assign n17845 = ~n16726 & n17844 ;
  assign n17846 = n17845 ^ n17480 ;
  assign n17847 = n17846 ^ n15997 ;
  assign n18106 = n17964 ^ n17847 ;
  assign n18107 = n18106 ^ x284 ;
  assign n18108 = n18107 ^ n18102 ;
  assign n18109 = n18108 ^ n18106 ;
  assign n18110 = ~n18105 & n18109 ;
  assign n18111 = n18110 ^ n18107 ;
  assign n17965 = n17964 ^ n17846 ;
  assign n17966 = n17847 & ~n17965 ;
  assign n17967 = n17966 ^ n15997 ;
  assign n18112 = n17967 ^ n16018 ;
  assign n17973 = n17384 ^ n17383 ;
  assign n17969 = n17572 ^ n17480 ;
  assign n17968 = n17842 ^ n17572 ;
  assign n17970 = n17969 ^ n17968 ;
  assign n17971 = n17841 & n17970 ;
  assign n17972 = n17971 ^ n17969 ;
  assign n17974 = n17973 ^ n17972 ;
  assign n17975 = n17974 ^ n17572 ;
  assign n17976 = ~n16747 & n17975 ;
  assign n17977 = n17976 ^ n17572 ;
  assign n18113 = n18112 ^ n17977 ;
  assign n18115 = n18113 ^ x283 ;
  assign n18114 = n18113 ^ n18106 ;
  assign n18116 = n18115 ^ n18114 ;
  assign n18117 = ~n18111 & n18116 ;
  assign n18118 = n18117 ^ n18115 ;
  assign n17978 = n17977 ^ n17967 ;
  assign n17979 = n17977 ^ n16018 ;
  assign n17980 = n17978 & ~n17979 ;
  assign n17981 = n17980 ^ n16018 ;
  assign n18119 = n17981 ^ n16039 ;
  assign n17987 = n17387 ^ n17385 ;
  assign n17983 = n17684 ^ n17572 ;
  assign n17982 = n17973 ^ n17684 ;
  assign n17984 = n17983 ^ n17982 ;
  assign n17985 = ~n17972 & ~n17984 ;
  assign n17986 = n17985 ^ n17983 ;
  assign n17988 = n17987 ^ n17986 ;
  assign n17989 = n17988 ^ n17684 ;
  assign n17990 = n16768 & ~n17989 ;
  assign n17991 = n17990 ^ n17684 ;
  assign n18120 = n18119 ^ n17991 ;
  assign n18122 = n18120 ^ x282 ;
  assign n18121 = n18120 ^ n18113 ;
  assign n18123 = n18122 ^ n18121 ;
  assign n18124 = n18118 & ~n18123 ;
  assign n18125 = n18124 ^ n18122 ;
  assign n18126 = n18118 ^ x282 ;
  assign n18127 = n18111 ^ x283 ;
  assign n18161 = n18129 & ~n18160 ;
  assign n18162 = n18127 & n18161 ;
  assign n18163 = ~n18126 & n18162 ;
  assign n18166 = n18163 ^ n18120 ;
  assign n18167 = n18125 & n18166 ;
  assign n18164 = n18163 ^ n18125 ;
  assign n18165 = x281 & n18164 ;
  assign n18168 = n18167 ^ n18165 ;
  assign n18002 = n17987 ^ n17684 ;
  assign n18003 = ~n17986 & ~n18002 ;
  assign n17999 = n17746 ^ n17388 ;
  assign n18000 = n17999 ^ n17389 ;
  assign n18001 = n18000 ^ n17987 ;
  assign n18004 = n18003 ^ n18001 ;
  assign n18005 = n18004 ^ n17746 ;
  assign n18006 = n16839 & ~n18005 ;
  assign n17996 = n17746 ^ n16127 ;
  assign n17995 = n16039 ^ x280 ;
  assign n17997 = n17996 ^ n17995 ;
  assign n17992 = n17991 ^ n17981 ;
  assign n17993 = n17991 ^ n16039 ;
  assign n17994 = n17992 & ~n17993 ;
  assign n17998 = n17997 ^ n17994 ;
  assign n18007 = n18006 ^ n17998 ;
  assign n18169 = n18168 ^ n18007 ;
  assign n17788 = n17787 ^ n17077 ;
  assign n18170 = n18169 ^ n17788 ;
  assign n18174 = n18162 ^ n18126 ;
  assign n18173 = n17775 ^ n17059 ;
  assign n18175 = n18174 ^ n18173 ;
  assign n18274 = n18273 ^ n18272 ;
  assign n18275 = n18273 ^ n17879 ;
  assign n18276 = n18274 & ~n18275 ;
  assign n18277 = n18276 ^ n17879 ;
  assign n18176 = n18161 ^ n18127 ;
  assign n18278 = n18277 ^ n18176 ;
  assign n18279 = n18174 ^ n17858 ;
  assign n18280 = n18279 ^ n18176 ;
  assign n18281 = n18280 ^ n18174 ;
  assign n18282 = ~n18278 & n18281 ;
  assign n18283 = n18282 ^ n18279 ;
  assign n18284 = ~n18175 & ~n18283 ;
  assign n18285 = n18284 ^ n18174 ;
  assign n18171 = n18125 ^ x281 ;
  assign n18172 = n18171 ^ n18163 ;
  assign n18286 = n18285 ^ n18172 ;
  assign n18287 = n18285 ^ n17897 ;
  assign n18288 = n18286 & ~n18287 ;
  assign n18289 = n18288 ^ n17897 ;
  assign n18290 = n18289 ^ n17788 ;
  assign n18291 = n18170 & ~n18290 ;
  assign n18292 = n18291 ^ n18169 ;
  assign n18293 = n18292 ^ n17911 ;
  assign n18294 = n17853 ^ n17701 ;
  assign n18295 = n18294 ^ n17853 ;
  assign n18296 = n18295 ^ n18292 ;
  assign n18297 = n18293 & ~n18296 ;
  assign n18298 = n18297 ^ n18294 ;
  assign n18443 = n17923 ^ n17853 ;
  assign n18299 = n17703 ^ n17701 ;
  assign n18442 = n18299 ^ n17923 ;
  assign n18444 = n18443 ^ n18442 ;
  assign n18445 = n18298 & ~n18444 ;
  assign n18446 = n18445 ^ n18443 ;
  assign n18457 = n17931 ^ n17923 ;
  assign n18447 = n17705 ^ n17704 ;
  assign n18456 = n18447 ^ n17931 ;
  assign n18458 = n18457 ^ n18456 ;
  assign n18459 = n18446 & n18458 ;
  assign n18460 = n18459 ^ n18457 ;
  assign n18461 = n17707 ^ n17706 ;
  assign n18468 = n18461 ^ n17931 ;
  assign n18469 = n18460 & ~n18468 ;
  assign n18470 = n18469 ^ n17931 ;
  assign n18467 = n17709 ^ n17708 ;
  assign n18471 = n18470 ^ n18467 ;
  assign n18627 = n18470 ^ n17848 ;
  assign n18628 = ~n18471 & ~n18627 ;
  assign n18629 = n18628 ^ n17848 ;
  assign n18647 = n18646 ^ n18629 ;
  assign n18630 = n17711 ^ n17710 ;
  assign n18648 = n18646 ^ n18630 ;
  assign n18649 = ~n18647 & n18648 ;
  assign n18645 = n18630 ^ n17949 ;
  assign n18650 = n18649 ^ n18645 ;
  assign n18668 = n17957 ^ n17949 ;
  assign n18651 = n17713 ^ n17712 ;
  assign n18667 = n18651 ^ n17957 ;
  assign n18669 = n18668 ^ n18667 ;
  assign n18670 = ~n18650 & ~n18669 ;
  assign n18671 = n18670 ^ n18668 ;
  assign n18751 = n17957 ^ n17843 ;
  assign n18672 = n17715 ^ n17714 ;
  assign n18750 = n18672 ^ n17843 ;
  assign n18752 = n18751 ^ n18750 ;
  assign n18753 = ~n18671 & ~n18752 ;
  assign n18754 = n18753 ^ n18751 ;
  assign n18788 = n17719 ^ n17718 ;
  assign n18790 = n18788 ^ n17843 ;
  assign n18755 = n17717 ^ n17716 ;
  assign n18789 = n18788 ^ n18755 ;
  assign n18791 = n18790 ^ n18789 ;
  assign n18792 = n18754 & ~n18791 ;
  assign n18793 = n18792 ^ n18790 ;
  assign n18808 = n17988 ^ n17974 ;
  assign n18807 = n18788 ^ n17988 ;
  assign n18809 = n18808 ^ n18807 ;
  assign n18810 = ~n18793 & ~n18809 ;
  assign n18811 = n18810 ^ n18808 ;
  assign n18812 = n17721 ^ n17720 ;
  assign n18841 = n18812 ^ n17988 ;
  assign n18842 = ~n18811 & ~n18841 ;
  assign n18839 = n17723 ^ n17722 ;
  assign n18840 = n18839 ^ n17988 ;
  assign n18843 = n18842 ^ n18840 ;
  assign n18844 = ~n17746 & n18843 ;
  assign n18836 = n18004 ^ n16839 ;
  assign n18835 = n16768 ^ x440 ;
  assign n18837 = n18836 ^ n18835 ;
  assign n18813 = n18812 ^ n18811 ;
  assign n18814 = n18813 ^ n17988 ;
  assign n18815 = ~n17684 & n18814 ;
  assign n18816 = n18815 ^ n17988 ;
  assign n18794 = ~n17572 & n18793 ;
  assign n18795 = n18794 ^ n17974 ;
  assign n18756 = n18755 ^ n18754 ;
  assign n18757 = n18756 ^ n17843 ;
  assign n18758 = n17480 & ~n18757 ;
  assign n18759 = n18758 ^ n17843 ;
  assign n18673 = n18672 ^ n18671 ;
  assign n18674 = n18673 ^ n17957 ;
  assign n18675 = n17341 & n18674 ;
  assign n18676 = n18675 ^ n17957 ;
  assign n18652 = n18651 ^ n18650 ;
  assign n18653 = n18652 ^ n17949 ;
  assign n18654 = n17320 & n18653 ;
  assign n18655 = n18654 ^ n17949 ;
  assign n18631 = n18630 ^ n18629 ;
  assign n18632 = ~n17825 & ~n18631 ;
  assign n18633 = n18632 ^ n17824 ;
  assign n18462 = n18461 ^ n18460 ;
  assign n18463 = n18462 ^ n17931 ;
  assign n18464 = ~n17129 & ~n18463 ;
  assign n18465 = n18464 ^ n17931 ;
  assign n18448 = n18447 ^ n18446 ;
  assign n18449 = n18448 ^ n17923 ;
  assign n18450 = ~n17116 & n18449 ;
  assign n18451 = n18450 ^ n17923 ;
  assign n18300 = n18299 ^ n18298 ;
  assign n18301 = n18300 ^ n17853 ;
  assign n18302 = ~n17103 & ~n18301 ;
  assign n18303 = n18302 ^ n17853 ;
  assign n18304 = n18303 ^ n16434 ;
  assign n18432 = n18292 ^ n17701 ;
  assign n18433 = ~n17090 & ~n18432 ;
  assign n18434 = n18433 ^ n17911 ;
  assign n18425 = n18289 ^ n18169 ;
  assign n18426 = n17077 & ~n18425 ;
  assign n18427 = n18426 ^ n17787 ;
  assign n18305 = ~n17059 & n18283 ;
  assign n18306 = n18305 ^ n17775 ;
  assign n18307 = n18306 ^ n16385 ;
  assign n18410 = n17047 & n18278 ;
  assign n18374 = n18373 ^ n18369 ;
  assign n18375 = ~n18370 & ~n18374 ;
  assign n18376 = n18375 ^ n16196 ;
  assign n18377 = n18376 ^ n16402 ;
  assign n18378 = ~n16954 & ~n18256 ;
  assign n18379 = n18378 ^ n18258 ;
  assign n18380 = n18379 ^ n18376 ;
  assign n18381 = n18377 & ~n18380 ;
  assign n18382 = n18381 ^ n16402 ;
  assign n18383 = n18382 ^ n16400 ;
  assign n18384 = n18261 ^ n18183 ;
  assign n18385 = n16949 & n18384 ;
  assign n18386 = n18385 ^ n18182 ;
  assign n18387 = n18386 ^ n18382 ;
  assign n18388 = n18383 & n18387 ;
  assign n18389 = n18388 ^ n16400 ;
  assign n18390 = n18389 ^ n16398 ;
  assign n18391 = ~n16944 & ~n18265 ;
  assign n18392 = n18391 ^ n18266 ;
  assign n18393 = n18392 ^ n18389 ;
  assign n18394 = ~n18390 & n18393 ;
  assign n18395 = n18394 ^ n16398 ;
  assign n18396 = n18395 ^ n16395 ;
  assign n18397 = n18269 ^ n18178 ;
  assign n18398 = ~n16939 & n18397 ;
  assign n18399 = n18398 ^ n18177 ;
  assign n18400 = n18399 ^ n18395 ;
  assign n18401 = n18396 & n18400 ;
  assign n18402 = n18401 ^ n16395 ;
  assign n18403 = n18402 ^ n16396 ;
  assign n18404 = ~n17042 & ~n18274 ;
  assign n18405 = n18404 ^ n17879 ;
  assign n18406 = n18405 ^ n18402 ;
  assign n18407 = n18403 & ~n18406 ;
  assign n18408 = n18407 ^ n16396 ;
  assign n18409 = n18408 ^ n17858 ;
  assign n18411 = n18410 ^ n18409 ;
  assign n18412 = n18306 ^ n16919 ;
  assign n18413 = n18412 ^ n18408 ;
  assign n18414 = n18413 ^ n18306 ;
  assign n18415 = ~n18411 & n18414 ;
  assign n18416 = n18415 ^ n18412 ;
  assign n18417 = n18307 & n18416 ;
  assign n18418 = n18417 ^ n16385 ;
  assign n18419 = n18418 ^ n16391 ;
  assign n18420 = n16934 & ~n18286 ;
  assign n18421 = n18420 ^ n17897 ;
  assign n18422 = n18421 ^ n18418 ;
  assign n18423 = n18419 & n18422 ;
  assign n18424 = n18423 ^ n16391 ;
  assign n18428 = n18427 ^ n18424 ;
  assign n18429 = n18427 ^ n16444 ;
  assign n18430 = n18428 & n18429 ;
  assign n18431 = n18430 ^ n16444 ;
  assign n18435 = n18434 ^ n18431 ;
  assign n18436 = n18434 ^ n16439 ;
  assign n18437 = n18435 & ~n18436 ;
  assign n18438 = n18437 ^ n16439 ;
  assign n18439 = n18438 ^ n18303 ;
  assign n18440 = ~n18304 & n18439 ;
  assign n18441 = n18440 ^ n16434 ;
  assign n18452 = n18451 ^ n18441 ;
  assign n18453 = n18451 ^ n16429 ;
  assign n18454 = n18452 & ~n18453 ;
  assign n18455 = n18454 ^ n16429 ;
  assign n18466 = n18465 ^ n18455 ;
  assign n18480 = n18455 ^ n16536 ;
  assign n18477 = n18466 & n18480 ;
  assign n18472 = ~n17791 & n18471 ;
  assign n18473 = n18472 ^ n17848 ;
  assign n18474 = n18473 ^ n16536 ;
  assign n18478 = n18477 ^ n18474 ;
  assign n18623 = n18473 ^ n16645 ;
  assign n18624 = ~n18478 & ~n18623 ;
  assign n18625 = n18624 ^ n16645 ;
  assign n18640 = n18633 ^ n18625 ;
  assign n18641 = n18633 ^ n17314 ;
  assign n18642 = ~n18640 & n18641 ;
  assign n18643 = n18642 ^ n17314 ;
  assign n18662 = n18655 ^ n18643 ;
  assign n18663 = n18655 ^ n16684 ;
  assign n18664 = ~n18662 & n18663 ;
  assign n18665 = n18664 ^ n16684 ;
  assign n18745 = n18676 ^ n18665 ;
  assign n18746 = n18676 ^ n16705 ;
  assign n18747 = n18745 & n18746 ;
  assign n18748 = n18747 ^ n16705 ;
  assign n18783 = n18759 ^ n18748 ;
  assign n18784 = n18759 ^ n16726 ;
  assign n18785 = ~n18783 & ~n18784 ;
  assign n18786 = n18785 ^ n16726 ;
  assign n18802 = n18795 ^ n18786 ;
  assign n18803 = n18795 ^ n16747 ;
  assign n18804 = ~n18802 & n18803 ;
  assign n18805 = n18804 ^ n16747 ;
  assign n18832 = n18816 ^ n18805 ;
  assign n18833 = n18816 ^ n16768 ;
  assign n18834 = n18832 & n18833 ;
  assign n18838 = n18837 ^ n18834 ;
  assign n18845 = n18844 ^ n18838 ;
  assign n18481 = n18480 ^ n18465 ;
  assign n18482 = n18481 ^ x432 ;
  assign n18485 = n18431 ^ n16439 ;
  assign n18486 = n18485 ^ n18434 ;
  assign n18487 = n18486 ^ x435 ;
  assign n18489 = n18405 ^ n18403 ;
  assign n18490 = n18489 ^ x424 ;
  assign n18549 = n18379 ^ n18377 ;
  assign n18551 = n18549 ^ x429 ;
  assign n18550 = n18549 ^ n18543 ;
  assign n18552 = n18551 ^ n18550 ;
  assign n18553 = n18548 & ~n18552 ;
  assign n18554 = n18553 ^ n18551 ;
  assign n18555 = n18386 ^ n18383 ;
  assign n18557 = n18555 ^ x428 ;
  assign n18556 = n18555 ^ n18549 ;
  assign n18558 = n18557 ^ n18556 ;
  assign n18559 = n18554 & ~n18558 ;
  assign n18560 = n18559 ^ n18557 ;
  assign n18561 = n18392 ^ n18390 ;
  assign n18563 = n18561 ^ x427 ;
  assign n18562 = n18561 ^ n18555 ;
  assign n18564 = n18563 ^ n18562 ;
  assign n18565 = ~n18560 & n18564 ;
  assign n18566 = n18565 ^ n18563 ;
  assign n18567 = n18399 ^ n18396 ;
  assign n18569 = n18567 ^ x426 ;
  assign n18568 = n18567 ^ n18561 ;
  assign n18570 = n18569 ^ n18568 ;
  assign n18571 = n18566 & ~n18570 ;
  assign n18572 = n18571 ^ n18569 ;
  assign n18574 = n18489 ^ x425 ;
  assign n18573 = n18567 ^ n18489 ;
  assign n18575 = n18574 ^ n18573 ;
  assign n18576 = n18572 & ~n18575 ;
  assign n18577 = n18576 ^ n18574 ;
  assign n18578 = n18490 & ~n18577 ;
  assign n18579 = n18578 ^ x424 ;
  assign n18488 = n18411 ^ n16919 ;
  assign n18580 = n18579 ^ n18488 ;
  assign n18581 = n18416 ^ n16385 ;
  assign n18582 = n18581 ^ x439 ;
  assign n18583 = n18582 ^ n18488 ;
  assign n18584 = n18583 ^ n18581 ;
  assign n18585 = ~n18580 & n18584 ;
  assign n18586 = n18585 ^ n18582 ;
  assign n18587 = n18421 ^ n18419 ;
  assign n18589 = n18587 ^ x438 ;
  assign n18588 = n18587 ^ n18581 ;
  assign n18590 = n18589 ^ n18588 ;
  assign n18591 = ~n18586 & n18590 ;
  assign n18592 = n18591 ^ n18589 ;
  assign n18593 = n18424 ^ n16444 ;
  assign n18594 = n18593 ^ n18427 ;
  assign n18596 = n18594 ^ x437 ;
  assign n18595 = n18594 ^ n18587 ;
  assign n18597 = n18596 ^ n18595 ;
  assign n18598 = ~n18592 & n18597 ;
  assign n18599 = n18598 ^ n18596 ;
  assign n18601 = n18486 ^ x436 ;
  assign n18600 = n18594 ^ n18486 ;
  assign n18602 = n18601 ^ n18600 ;
  assign n18603 = n18599 & ~n18602 ;
  assign n18604 = n18603 ^ n18601 ;
  assign n18605 = ~n18487 & n18604 ;
  assign n18606 = n18605 ^ x435 ;
  assign n18483 = n18438 ^ n16434 ;
  assign n18484 = n18483 ^ n18303 ;
  assign n18607 = n18606 ^ n18484 ;
  assign n18608 = n18441 ^ n16429 ;
  assign n18609 = n18608 ^ n18451 ;
  assign n18610 = n18609 ^ x434 ;
  assign n18611 = n18610 ^ n18606 ;
  assign n18612 = n18611 ^ n18609 ;
  assign n18613 = n18607 & n18612 ;
  assign n18614 = n18613 ^ n18610 ;
  assign n18616 = n18481 ^ x433 ;
  assign n18615 = n18609 ^ n18481 ;
  assign n18617 = n18616 ^ n18615 ;
  assign n18618 = n18614 & ~n18617 ;
  assign n18619 = n18618 ^ n18616 ;
  assign n18620 = ~n18482 & n18619 ;
  assign n18621 = n18620 ^ x432 ;
  assign n18479 = n18478 ^ n16645 ;
  assign n18622 = n18621 ^ n18479 ;
  assign n18626 = n18625 ^ n17314 ;
  assign n18634 = n18633 ^ n18626 ;
  assign n18635 = n18634 ^ x447 ;
  assign n18636 = n18635 ^ n18479 ;
  assign n18637 = n18636 ^ n18634 ;
  assign n18638 = n18622 & ~n18637 ;
  assign n18639 = n18638 ^ n18635 ;
  assign n18644 = n18643 ^ n16684 ;
  assign n18656 = n18655 ^ n18644 ;
  assign n18658 = n18656 ^ x446 ;
  assign n18657 = n18656 ^ n18634 ;
  assign n18659 = n18658 ^ n18657 ;
  assign n18660 = n18639 & ~n18659 ;
  assign n18661 = n18660 ^ n18658 ;
  assign n18666 = n18665 ^ n16705 ;
  assign n18677 = n18676 ^ n18666 ;
  assign n18679 = n18677 ^ x445 ;
  assign n18678 = n18677 ^ n18656 ;
  assign n18680 = n18679 ^ n18678 ;
  assign n18681 = n18661 & ~n18680 ;
  assign n18682 = n18681 ^ n18679 ;
  assign n18749 = n18748 ^ n16726 ;
  assign n18760 = n18759 ^ n18749 ;
  assign n18762 = n18760 ^ x444 ;
  assign n18761 = n18760 ^ n18677 ;
  assign n18763 = n18762 ^ n18761 ;
  assign n18764 = n18682 & ~n18763 ;
  assign n18765 = n18764 ^ n18762 ;
  assign n18787 = n18786 ^ n16747 ;
  assign n18796 = n18795 ^ n18787 ;
  assign n18798 = n18796 ^ x443 ;
  assign n18797 = n18796 ^ n18760 ;
  assign n18799 = n18798 ^ n18797 ;
  assign n18800 = n18765 & ~n18799 ;
  assign n18801 = n18800 ^ n18798 ;
  assign n18806 = n18805 ^ n16768 ;
  assign n18817 = n18816 ^ n18806 ;
  assign n18819 = n18817 ^ x442 ;
  assign n18818 = n18817 ^ n18796 ;
  assign n18820 = n18819 ^ n18818 ;
  assign n18821 = n18801 & ~n18820 ;
  assign n18822 = n18821 ^ n18819 ;
  assign n18766 = n18765 ^ x443 ;
  assign n18683 = n18682 ^ x444 ;
  assign n18705 = n18703 & ~n18704 ;
  assign n18706 = n18554 ^ x428 ;
  assign n18707 = ~n18705 & n18706 ;
  assign n18708 = n18560 ^ x427 ;
  assign n18709 = ~n18707 & n18708 ;
  assign n18710 = n18566 ^ x426 ;
  assign n18711 = ~n18709 & n18710 ;
  assign n18712 = n18572 ^ x425 ;
  assign n18713 = n18711 & n18712 ;
  assign n18714 = n18577 ^ x424 ;
  assign n18715 = n18713 & ~n18714 ;
  assign n18716 = n18579 ^ x439 ;
  assign n18717 = n18716 ^ n18488 ;
  assign n18718 = n18715 & ~n18717 ;
  assign n18719 = n18586 ^ x438 ;
  assign n18720 = n18718 & ~n18719 ;
  assign n18721 = n18592 ^ x437 ;
  assign n18722 = ~n18720 & n18721 ;
  assign n18723 = n18599 ^ x436 ;
  assign n18724 = n18722 & ~n18723 ;
  assign n18725 = n18604 ^ x435 ;
  assign n18726 = n18724 & ~n18725 ;
  assign n18727 = n18607 ^ x434 ;
  assign n18728 = ~n18726 & n18727 ;
  assign n18729 = n18614 ^ x433 ;
  assign n18730 = n18728 & n18729 ;
  assign n18731 = n18619 ^ x432 ;
  assign n18732 = n18730 & n18731 ;
  assign n18733 = n18621 ^ x447 ;
  assign n18734 = n18733 ^ n18479 ;
  assign n18735 = n18732 & n18734 ;
  assign n18736 = n18639 ^ x446 ;
  assign n18737 = ~n18735 & ~n18736 ;
  assign n18738 = n18661 ^ x445 ;
  assign n18739 = n18737 & ~n18738 ;
  assign n18767 = n18683 & ~n18739 ;
  assign n18824 = ~n18766 & ~n18767 ;
  assign n18825 = n18801 ^ x442 ;
  assign n18826 = ~n18824 & n18825 ;
  assign n18827 = n18826 ^ n18817 ;
  assign n18830 = n18822 & ~n18827 ;
  assign n18823 = n18822 ^ n18817 ;
  assign n18828 = n18827 ^ n18823 ;
  assign n18829 = ~x441 & n18828 ;
  assign n18831 = n18830 ^ n18829 ;
  assign n18846 = n18845 ^ n18831 ;
  assign n18781 = n18231 ^ n18209 ;
  assign n18782 = n18781 ^ n18207 ;
  assign n18847 = n18846 ^ n18782 ;
  assign n18850 = n18229 ^ n18213 ;
  assign n18848 = n18822 ^ x441 ;
  assign n18849 = n18848 ^ n18826 ;
  assign n18851 = n18850 ^ n18849 ;
  assign n18854 = n18825 ^ n18824 ;
  assign n18852 = n18225 ^ n18217 ;
  assign n18853 = n18852 ^ n18215 ;
  assign n18855 = n18854 ^ n18853 ;
  assign n17727 = n17726 ^ n17725 ;
  assign n18740 = n18739 ^ n18683 ;
  assign n18743 = n17727 & n18740 ;
  assign n18742 = n18222 ^ n18221 ;
  assign n18744 = n18743 ^ n18742 ;
  assign n18768 = n18767 ^ n18766 ;
  assign n18856 = n18768 ^ n18743 ;
  assign n18857 = ~n18744 & n18856 ;
  assign n18858 = n18857 ^ n18768 ;
  assign n18859 = n18858 ^ n18853 ;
  assign n18860 = ~n18855 & n18859 ;
  assign n18861 = n18860 ^ n18854 ;
  assign n18862 = n18861 ^ n18849 ;
  assign n18863 = n18851 & ~n18862 ;
  assign n18864 = n18863 ^ n18850 ;
  assign n18865 = n18864 ^ n18782 ;
  assign n18866 = n18847 & ~n18865 ;
  assign n18867 = n18866 ^ n18846 ;
  assign n18869 = n18868 ^ n18867 ;
  assign n18870 = n18238 ^ n18201 ;
  assign n18871 = n18870 ^ n18686 ;
  assign n18872 = n18871 ^ n18870 ;
  assign n18873 = n18872 ^ n18867 ;
  assign n18874 = n18869 & ~n18873 ;
  assign n18875 = n18874 ^ n18871 ;
  assign n18877 = n18241 ^ n18197 ;
  assign n18879 = n18877 ^ n18870 ;
  assign n18876 = n18687 ^ n18686 ;
  assign n18878 = n18877 ^ n18876 ;
  assign n18880 = n18879 ^ n18878 ;
  assign n18881 = ~n18875 & ~n18880 ;
  assign n18882 = n18881 ^ n18879 ;
  assign n18885 = n18877 ^ n18777 ;
  assign n18883 = n18689 ^ n18688 ;
  assign n18884 = n18883 ^ n18777 ;
  assign n18886 = n18885 ^ n18884 ;
  assign n18887 = ~n18882 & n18886 ;
  assign n18888 = n18887 ^ n18885 ;
  assign n18889 = n18780 & n18888 ;
  assign n18778 = n18777 ^ n18774 ;
  assign n18890 = n18889 ^ n18778 ;
  assign n18891 = n18775 & n18890 ;
  assign n18772 = n18695 ^ n18694 ;
  assign n18773 = n18772 ^ n18771 ;
  assign n18892 = n18891 ^ n18773 ;
  assign n18896 = n18253 ^ n18188 ;
  assign n18893 = n18258 ^ n18255 ;
  assign n18894 = n18893 ^ n18185 ;
  assign n18897 = n18896 ^ n18894 ;
  assign n18895 = n18894 ^ n18772 ;
  assign n18898 = n18897 ^ n18895 ;
  assign n18899 = n18892 & n18898 ;
  assign n18900 = n18899 ^ n18895 ;
  assign n18901 = n18696 ^ n18684 ;
  assign n18948 = n18901 ^ n18894 ;
  assign n18949 = n18900 & ~n18948 ;
  assign n18950 = n18949 ^ n18894 ;
  assign n18947 = n18698 ^ n18697 ;
  assign n18951 = n18950 ^ n18947 ;
  assign n18955 = n18262 ^ n18183 ;
  assign n18952 = n18266 ^ n18264 ;
  assign n18953 = n18952 ^ n18180 ;
  assign n18954 = n18953 ^ n18950 ;
  assign n18956 = n18955 ^ n18954 ;
  assign n18957 = n18956 ^ n18953 ;
  assign n18958 = ~n18951 & n18957 ;
  assign n18959 = n18958 ^ n18954 ;
  assign n18962 = n18953 ^ n18770 ;
  assign n18960 = n18700 ^ n18699 ;
  assign n18961 = n18960 ^ n18770 ;
  assign n18963 = n18962 ^ n18961 ;
  assign n18964 = ~n18959 & n18963 ;
  assign n18965 = n18964 ^ n18962 ;
  assign n18966 = n18702 ^ n18701 ;
  assign n18967 = n18966 ^ n18770 ;
  assign n18968 = n18965 & ~n18967 ;
  assign n18972 = n18971 ^ n18968 ;
  assign n19130 = n18973 ^ n18972 ;
  assign n19131 = n19130 ^ n18970 ;
  assign n19132 = n17879 & n19131 ;
  assign n19133 = n19132 ^ n18970 ;
  assign n19070 = n18883 ^ n18882 ;
  assign n19071 = n19070 ^ n18877 ;
  assign n19072 = ~n18196 & ~n19071 ;
  assign n19073 = n19072 ^ n18877 ;
  assign n19048 = n18864 ^ n18846 ;
  assign n19049 = n18209 & n19048 ;
  assign n19050 = n19049 ^ n18782 ;
  assign n19042 = n18212 & n18862 ;
  assign n19043 = n19042 ^ n18850 ;
  assign n18917 = n18858 ^ n18854 ;
  assign n18918 = ~n18217 & n18917 ;
  assign n18919 = n18918 ^ n18853 ;
  assign n18905 = ~n17726 & ~n18740 ;
  assign n18906 = n18905 ^ n17725 ;
  assign n18907 = n17436 & ~n18906 ;
  assign n18908 = n18907 ^ n17439 ;
  assign n18903 = ~n18220 & n18856 ;
  assign n18904 = n18903 ^ n18742 ;
  assign n18913 = n18907 ^ n18904 ;
  assign n18914 = ~n18908 & ~n18913 ;
  assign n18915 = n18914 ^ n17439 ;
  assign n19038 = n18919 ^ n18915 ;
  assign n19039 = n18919 ^ n17434 ;
  assign n19040 = ~n19038 & ~n19039 ;
  assign n19041 = n19040 ^ n17434 ;
  assign n19044 = n19043 ^ n19041 ;
  assign n19045 = n19043 ^ n17431 ;
  assign n19046 = ~n19044 & ~n19045 ;
  assign n19047 = n19046 ^ n17431 ;
  assign n19051 = n19050 ^ n19047 ;
  assign n19052 = n19050 ^ n17427 ;
  assign n19053 = n19051 & n19052 ;
  assign n19054 = n19053 ^ n17427 ;
  assign n19055 = n19054 ^ n17424 ;
  assign n19056 = n18867 ^ n18686 ;
  assign n19057 = ~n18204 & ~n19056 ;
  assign n19058 = n19057 ^ n18868 ;
  assign n19059 = n19058 ^ n19054 ;
  assign n19060 = ~n19055 & n19059 ;
  assign n19061 = n19060 ^ n17424 ;
  assign n19062 = n19061 ^ n17420 ;
  assign n19063 = n18876 ^ n18875 ;
  assign n19064 = n19063 ^ n18870 ;
  assign n19065 = ~n18200 & n19064 ;
  assign n19066 = n19065 ^ n18870 ;
  assign n19067 = n19066 ^ n19061 ;
  assign n19068 = n19062 & n19067 ;
  assign n19069 = n19068 ^ n17420 ;
  assign n19074 = n19073 ^ n19069 ;
  assign n19075 = n19073 ^ n17416 ;
  assign n19076 = ~n19074 & ~n19075 ;
  assign n19077 = n19076 ^ n17416 ;
  assign n19078 = n19077 ^ n17412 ;
  assign n19079 = n18888 ^ n18779 ;
  assign n19080 = n19079 ^ n18777 ;
  assign n19081 = n18246 & n19080 ;
  assign n19082 = n19081 ^ n18777 ;
  assign n19083 = n19082 ^ n19077 ;
  assign n19084 = n19078 & n19083 ;
  assign n19085 = n19084 ^ n17412 ;
  assign n19086 = n19085 ^ n17015 ;
  assign n19087 = n18890 ^ n18771 ;
  assign n19088 = n19087 ^ n18774 ;
  assign n19089 = ~n18191 & ~n19088 ;
  assign n19090 = n19089 ^ n18774 ;
  assign n19091 = n19090 ^ n19085 ;
  assign n19092 = ~n19086 & ~n19091 ;
  assign n19093 = n19092 ^ n17015 ;
  assign n19094 = n19093 ^ n17022 ;
  assign n19095 = n18187 & n18892 ;
  assign n19096 = n19095 ^ n18896 ;
  assign n19097 = n19096 ^ n19093 ;
  assign n19098 = n19094 & n19097 ;
  assign n19099 = n19098 ^ n17022 ;
  assign n19100 = n19099 ^ n16954 ;
  assign n18902 = n18901 ^ n18900 ;
  assign n19101 = n18902 ^ n18894 ;
  assign n19102 = ~n18258 & ~n19101 ;
  assign n19103 = n19102 ^ n18894 ;
  assign n19104 = n19103 ^ n19099 ;
  assign n19105 = n19100 & n19104 ;
  assign n19106 = n19105 ^ n16954 ;
  assign n19107 = n19106 ^ n16949 ;
  assign n19108 = n18182 & ~n18951 ;
  assign n19109 = n19108 ^ n18955 ;
  assign n19110 = n19109 ^ n19106 ;
  assign n19111 = ~n19107 & n19110 ;
  assign n19112 = n19111 ^ n16949 ;
  assign n19113 = n19112 ^ n16944 ;
  assign n19114 = n18960 ^ n18959 ;
  assign n19115 = n19114 ^ n18953 ;
  assign n19116 = n18266 & ~n19115 ;
  assign n19117 = n19116 ^ n18953 ;
  assign n19118 = n19117 ^ n19112 ;
  assign n19119 = ~n19113 & n19118 ;
  assign n19120 = n19119 ^ n16944 ;
  assign n19121 = n19120 ^ n16939 ;
  assign n19122 = n18966 ^ n18965 ;
  assign n19123 = n19122 ^ n18770 ;
  assign n19124 = ~n18177 & ~n19123 ;
  assign n19125 = n19124 ^ n18770 ;
  assign n19126 = n19125 ^ n19120 ;
  assign n19127 = n19121 & ~n19126 ;
  assign n19128 = n19127 ^ n16939 ;
  assign n19129 = n19128 ^ n17042 ;
  assign n19287 = n19133 ^ n19129 ;
  assign n19288 = n19287 ^ x72 ;
  assign n18910 = n18906 ^ n17436 ;
  assign n18911 = x71 & ~n18910 ;
  assign n18909 = n18908 ^ n18904 ;
  assign n18912 = n18911 ^ n18909 ;
  assign n18916 = n18915 ^ n17434 ;
  assign n18920 = n18919 ^ n18916 ;
  assign n18921 = n18920 ^ x70 ;
  assign n18922 = n18921 ^ n18909 ;
  assign n18923 = n18922 ^ n18920 ;
  assign n18924 = n18912 & ~n18923 ;
  assign n18925 = n18924 ^ n18921 ;
  assign n19289 = n19041 ^ n17431 ;
  assign n19290 = n19289 ^ n19043 ;
  assign n19292 = n19290 ^ x69 ;
  assign n19291 = n19290 ^ n18920 ;
  assign n19293 = n19292 ^ n19291 ;
  assign n19294 = ~n18925 & n19293 ;
  assign n19295 = n19294 ^ n19292 ;
  assign n19296 = n19047 ^ n17427 ;
  assign n19297 = n19296 ^ n19050 ;
  assign n19299 = n19297 ^ x68 ;
  assign n19298 = n19297 ^ n19290 ;
  assign n19300 = n19299 ^ n19298 ;
  assign n19301 = n19295 & ~n19300 ;
  assign n19302 = n19301 ^ n19299 ;
  assign n19303 = n19058 ^ n19055 ;
  assign n19305 = n19303 ^ x67 ;
  assign n19304 = n19303 ^ n19297 ;
  assign n19306 = n19305 ^ n19304 ;
  assign n19307 = n19302 & ~n19306 ;
  assign n19308 = n19307 ^ n19305 ;
  assign n19309 = n19066 ^ n19062 ;
  assign n19311 = n19309 ^ x66 ;
  assign n19310 = n19309 ^ n19303 ;
  assign n19312 = n19311 ^ n19310 ;
  assign n19313 = ~n19308 & n19312 ;
  assign n19314 = n19313 ^ n19311 ;
  assign n19315 = n19069 ^ n17416 ;
  assign n19316 = n19315 ^ n19073 ;
  assign n19318 = n19316 ^ x65 ;
  assign n19317 = n19316 ^ n19309 ;
  assign n19319 = n19318 ^ n19317 ;
  assign n19320 = ~n19314 & n19319 ;
  assign n19321 = n19320 ^ n19318 ;
  assign n19322 = n19082 ^ n19078 ;
  assign n19324 = n19322 ^ x64 ;
  assign n19323 = n19322 ^ n19316 ;
  assign n19325 = n19324 ^ n19323 ;
  assign n19326 = ~n19321 & n19325 ;
  assign n19327 = n19326 ^ n19324 ;
  assign n19328 = n19090 ^ n19086 ;
  assign n19330 = n19328 ^ x79 ;
  assign n19329 = n19328 ^ n19322 ;
  assign n19331 = n19330 ^ n19329 ;
  assign n19332 = n19327 & ~n19331 ;
  assign n19333 = n19332 ^ n19330 ;
  assign n19334 = n19096 ^ n19094 ;
  assign n19336 = n19334 ^ x78 ;
  assign n19335 = n19334 ^ n19328 ;
  assign n19337 = n19336 ^ n19335 ;
  assign n19338 = n19333 & ~n19337 ;
  assign n19339 = n19338 ^ n19336 ;
  assign n19340 = n19103 ^ n19100 ;
  assign n19342 = n19340 ^ x77 ;
  assign n19341 = n19340 ^ n19334 ;
  assign n19343 = n19342 ^ n19341 ;
  assign n19344 = ~n19339 & n19343 ;
  assign n19345 = n19344 ^ n19342 ;
  assign n19346 = n19109 ^ n19107 ;
  assign n19348 = n19346 ^ x76 ;
  assign n19347 = n19346 ^ n19340 ;
  assign n19349 = n19348 ^ n19347 ;
  assign n19350 = ~n19345 & n19349 ;
  assign n19351 = n19350 ^ n19348 ;
  assign n19352 = n19117 ^ n19113 ;
  assign n19354 = n19352 ^ x75 ;
  assign n19353 = n19352 ^ n19346 ;
  assign n19355 = n19354 ^ n19353 ;
  assign n19356 = n19351 & ~n19355 ;
  assign n19357 = n19356 ^ n19354 ;
  assign n19358 = n19125 ^ n19121 ;
  assign n19360 = n19358 ^ x74 ;
  assign n19359 = n19358 ^ n19352 ;
  assign n19361 = n19360 ^ n19359 ;
  assign n19362 = ~n19357 & n19361 ;
  assign n19363 = n19362 ^ n19360 ;
  assign n19365 = n19287 ^ x73 ;
  assign n19364 = n19358 ^ n19287 ;
  assign n19366 = n19365 ^ n19364 ;
  assign n19367 = n19363 & ~n19366 ;
  assign n19368 = n19367 ^ n19365 ;
  assign n19369 = ~n19288 & n19368 ;
  assign n19370 = n19369 ^ x72 ;
  assign n18974 = n18973 ^ n18970 ;
  assign n18975 = n18972 & n18974 ;
  assign n18976 = n18975 ^ n18970 ;
  assign n18946 = n18706 ^ n18705 ;
  assign n18977 = n18976 ^ n18946 ;
  assign n19137 = n17858 & ~n18977 ;
  assign n18978 = n18176 ^ n17858 ;
  assign n18979 = n18978 ^ n18277 ;
  assign n19138 = n19137 ^ n18979 ;
  assign n19285 = n19138 ^ n17047 ;
  assign n19134 = n19133 ^ n19128 ;
  assign n19135 = n19129 & ~n19134 ;
  assign n19136 = n19135 ^ n17042 ;
  assign n19286 = n19285 ^ n19136 ;
  assign n19371 = n19370 ^ n19286 ;
  assign n19139 = n19138 ^ n19136 ;
  assign n18983 = n18708 ^ n18707 ;
  assign n18980 = n18979 ^ n18946 ;
  assign n18981 = ~n18977 & ~n18980 ;
  assign n18982 = n18981 ^ n18976 ;
  assign n18984 = n18983 ^ n18982 ;
  assign n19035 = n18173 & ~n18984 ;
  assign n19036 = n19035 ^ n18283 ;
  assign n19140 = n19036 ^ n17047 ;
  assign n19141 = n19140 ^ n19136 ;
  assign n19142 = n19141 ^ n19036 ;
  assign n19143 = n19139 & ~n19142 ;
  assign n19144 = n19143 ^ n19140 ;
  assign n19372 = n19144 ^ n17059 ;
  assign n19373 = n19372 ^ x87 ;
  assign n19374 = n19373 ^ n19286 ;
  assign n19375 = n19374 ^ n19372 ;
  assign n19376 = n19371 & ~n19375 ;
  assign n19377 = n19376 ^ n19373 ;
  assign n18993 = n18710 ^ n18709 ;
  assign n18988 = n18287 ^ n18172 ;
  assign n18985 = n18283 ^ n18173 ;
  assign n18989 = n18988 ^ n18985 ;
  assign n18986 = n18985 ^ n18982 ;
  assign n18987 = ~n18984 & n18986 ;
  assign n18990 = n18989 ^ n18987 ;
  assign n19148 = n18993 ^ n18990 ;
  assign n19149 = n19148 ^ n18988 ;
  assign n19150 = n17897 & ~n19149 ;
  assign n19151 = n19150 ^ n18988 ;
  assign n19037 = n19036 ^ n17059 ;
  assign n19145 = n19037 & n19144 ;
  assign n19146 = n19145 ^ n17059 ;
  assign n19147 = n19146 ^ n16934 ;
  assign n19378 = n19151 ^ n19147 ;
  assign n19380 = n19378 ^ x86 ;
  assign n19379 = n19378 ^ n19372 ;
  assign n19381 = n19380 ^ n19379 ;
  assign n19382 = ~n19377 & n19381 ;
  assign n19383 = n19382 ^ n19380 ;
  assign n18998 = n18712 ^ n18711 ;
  assign n18991 = n18290 ^ n18169 ;
  assign n18992 = n18991 ^ n18988 ;
  assign n18994 = n18993 ^ n18992 ;
  assign n18995 = n18994 ^ n18991 ;
  assign n18996 = n18990 & ~n18995 ;
  assign n18997 = n18996 ^ n18992 ;
  assign n19156 = n18998 ^ n18997 ;
  assign n19157 = n19156 ^ n18991 ;
  assign n19158 = n17788 & n19157 ;
  assign n19159 = n19158 ^ n18991 ;
  assign n19152 = n19151 ^ n19146 ;
  assign n19153 = ~n19147 & ~n19152 ;
  assign n19154 = n19153 ^ n16934 ;
  assign n19155 = n19154 ^ n17077 ;
  assign n19384 = n19159 ^ n19155 ;
  assign n19386 = n19384 ^ x85 ;
  assign n19385 = n19384 ^ n19378 ;
  assign n19387 = n19386 ^ n19385 ;
  assign n19388 = ~n19383 & n19387 ;
  assign n19389 = n19388 ^ n19386 ;
  assign n18941 = n17911 ^ n17701 ;
  assign n18942 = n18941 ^ n18292 ;
  assign n19000 = n18991 ^ n18942 ;
  assign n18999 = n18998 ^ n18942 ;
  assign n19001 = n19000 ^ n18999 ;
  assign n19002 = ~n18997 & ~n19001 ;
  assign n19003 = n19002 ^ n19000 ;
  assign n18944 = n18714 ^ n18713 ;
  assign n19164 = n19003 ^ n18944 ;
  assign n19165 = n19164 ^ n18942 ;
  assign n19166 = ~n17911 & n19165 ;
  assign n19167 = n19166 ^ n18942 ;
  assign n19160 = n19159 ^ n19154 ;
  assign n19161 = n19155 & ~n19160 ;
  assign n19162 = n19161 ^ n17077 ;
  assign n19163 = n19162 ^ n17090 ;
  assign n19390 = n19167 ^ n19163 ;
  assign n19392 = n19390 ^ x84 ;
  assign n19391 = n19390 ^ n19384 ;
  assign n19393 = n19392 ^ n19391 ;
  assign n19394 = ~n19389 & n19393 ;
  assign n19395 = n19394 ^ n19392 ;
  assign n19008 = n18717 ^ n18715 ;
  assign n18945 = n18944 ^ n18942 ;
  assign n19004 = n18945 & n19003 ;
  assign n18943 = n18942 ^ n18300 ;
  assign n19005 = n19004 ^ n18943 ;
  assign n19172 = n19008 ^ n19005 ;
  assign n19173 = n19172 ^ n18300 ;
  assign n19174 = ~n17853 & n19173 ;
  assign n19175 = n19174 ^ n18300 ;
  assign n19168 = n19167 ^ n19162 ;
  assign n19169 = ~n19163 & ~n19168 ;
  assign n19170 = n19169 ^ n17090 ;
  assign n19171 = n19170 ^ n17103 ;
  assign n19396 = n19175 ^ n19171 ;
  assign n19398 = n19396 ^ x83 ;
  assign n19397 = n19396 ^ n19390 ;
  assign n19399 = n19398 ^ n19397 ;
  assign n19400 = n19395 & ~n19399 ;
  assign n19401 = n19400 ^ n19398 ;
  assign n19012 = n18719 ^ n18718 ;
  assign n19006 = n18448 ^ n18300 ;
  assign n19007 = n19006 ^ n18448 ;
  assign n19009 = n19008 ^ n19007 ;
  assign n19010 = n19005 & n19009 ;
  assign n19011 = n19010 ^ n19006 ;
  assign n19180 = n19012 ^ n19011 ;
  assign n19181 = n19180 ^ n18448 ;
  assign n19182 = ~n17923 & n19181 ;
  assign n19183 = n19182 ^ n18448 ;
  assign n19176 = n19175 ^ n19170 ;
  assign n19177 = n19171 & n19176 ;
  assign n19178 = n19177 ^ n17103 ;
  assign n19179 = n19178 ^ n17116 ;
  assign n19402 = n19183 ^ n19179 ;
  assign n19404 = n19402 ^ x82 ;
  assign n19403 = n19402 ^ n19396 ;
  assign n19405 = n19404 ^ n19403 ;
  assign n19406 = ~n19401 & n19405 ;
  assign n19407 = n19406 ^ n19404 ;
  assign n19184 = n19183 ^ n19178 ;
  assign n19185 = n19179 & ~n19184 ;
  assign n19186 = n19185 ^ n17116 ;
  assign n19282 = n19186 ^ n17129 ;
  assign n19014 = n18462 ^ n18448 ;
  assign n19013 = n19012 ^ n18462 ;
  assign n19015 = n19014 ^ n19013 ;
  assign n19016 = ~n19011 & ~n19015 ;
  assign n19017 = n19016 ^ n19014 ;
  assign n18939 = n18721 ^ n18720 ;
  assign n19187 = n19017 ^ n18939 ;
  assign n19188 = n19187 ^ n18462 ;
  assign n19189 = ~n17931 & n19188 ;
  assign n19190 = n19189 ^ n18462 ;
  assign n19283 = n19282 ^ n19190 ;
  assign n19409 = n19283 ^ x81 ;
  assign n19408 = n19402 ^ n19283 ;
  assign n19410 = n19409 ^ n19408 ;
  assign n19411 = n19407 & ~n19410 ;
  assign n19412 = n19411 ^ n19409 ;
  assign n19496 = n19412 ^ x80 ;
  assign n19456 = n19321 ^ x64 ;
  assign n19457 = n19295 ^ x68 ;
  assign n19458 = n19302 ^ x67 ;
  assign n19459 = n19457 & n19458 ;
  assign n19460 = n19308 ^ x66 ;
  assign n19461 = n19459 & ~n19460 ;
  assign n19462 = n19314 ^ x65 ;
  assign n19463 = n19461 & ~n19462 ;
  assign n19464 = ~n19456 & n19463 ;
  assign n19465 = n19327 ^ x79 ;
  assign n19466 = n19464 & n19465 ;
  assign n19467 = n19333 ^ x78 ;
  assign n19468 = n19466 & n19467 ;
  assign n19469 = n19339 ^ x77 ;
  assign n19470 = ~n19468 & n19469 ;
  assign n19471 = n19345 ^ x76 ;
  assign n19472 = n19470 & n19471 ;
  assign n19473 = n19351 ^ x75 ;
  assign n19474 = n19472 & ~n19473 ;
  assign n19475 = n19357 ^ x74 ;
  assign n19476 = ~n19474 & ~n19475 ;
  assign n19477 = n19363 ^ x73 ;
  assign n19478 = ~n19476 & ~n19477 ;
  assign n19479 = n19368 ^ x72 ;
  assign n19480 = ~n19478 & n19479 ;
  assign n19481 = n19370 ^ x87 ;
  assign n19482 = n19481 ^ n19286 ;
  assign n19483 = n19480 & n19482 ;
  assign n19484 = n19377 ^ x86 ;
  assign n19485 = n19483 & ~n19484 ;
  assign n19486 = n19383 ^ x85 ;
  assign n19487 = n19485 & ~n19486 ;
  assign n19488 = n19389 ^ x84 ;
  assign n19489 = n19487 & ~n19488 ;
  assign n19490 = n19395 ^ x83 ;
  assign n19491 = ~n19489 & ~n19490 ;
  assign n19492 = n19401 ^ x82 ;
  assign n19493 = ~n19491 & ~n19492 ;
  assign n19494 = n19407 ^ x81 ;
  assign n19495 = n19493 & n19494 ;
  assign n19536 = n19496 ^ n19495 ;
  assign n18741 = n18740 ^ n17727 ;
  assign n19923 = n19536 ^ n18741 ;
  assign n19633 = n17727 & ~n19536 ;
  assign n19634 = n19633 ^ n18740 ;
  assign n19707 = n19634 ^ n17726 ;
  assign n19882 = n19707 ^ x231 ;
  assign n19708 = x231 & ~n19707 ;
  assign n19883 = n19708 ^ x230 ;
  assign n19284 = n19283 ^ x80 ;
  assign n19413 = n19284 & ~n19412 ;
  assign n19414 = n19413 ^ x80 ;
  assign n19498 = n19414 ^ x95 ;
  assign n19191 = n19190 ^ n19186 ;
  assign n18940 = n18939 ^ n18462 ;
  assign n19018 = ~n18940 & ~n19017 ;
  assign n19019 = n19018 ^ n18462 ;
  assign n18938 = n18723 ^ n18722 ;
  assign n19020 = n19019 ^ n18938 ;
  assign n19192 = n17848 & ~n19020 ;
  assign n19021 = n18467 ^ n17848 ;
  assign n19022 = n19021 ^ n18470 ;
  assign n19193 = n19192 ^ n19022 ;
  assign n19194 = n19193 ^ n17129 ;
  assign n19195 = n19194 ^ n19186 ;
  assign n19196 = n19195 ^ n19193 ;
  assign n19197 = n19191 & n19196 ;
  assign n19198 = n19197 ^ n19194 ;
  assign n19281 = n19198 ^ n17791 ;
  assign n19499 = n19498 ^ n19281 ;
  assign n19497 = n19495 & ~n19496 ;
  assign n19539 = n19499 ^ n19497 ;
  assign n19537 = n18741 & n19536 ;
  assign n19540 = n19539 ^ n19537 ;
  assign n19637 = n18742 & ~n19540 ;
  assign n18769 = n18768 ^ n18744 ;
  assign n19638 = n19637 ^ n18769 ;
  assign n19635 = ~n17726 & n19634 ;
  assign n19636 = n19635 ^ n18220 ;
  assign n19706 = n19638 ^ n19636 ;
  assign n19884 = n19883 ^ n19706 ;
  assign n19885 = ~n19882 & ~n19884 ;
  assign n19709 = n19708 ^ n19706 ;
  assign n19639 = n19638 ^ n19635 ;
  assign n19640 = ~n19636 & ~n19639 ;
  assign n19641 = n19640 ^ n18220 ;
  assign n19710 = n19641 ^ n18217 ;
  assign n19538 = n19537 ^ n18769 ;
  assign n19541 = n19538 & n19540 ;
  assign n19542 = n19541 ^ n18769 ;
  assign n19415 = n19414 ^ n19281 ;
  assign n18934 = n18646 ^ n18631 ;
  assign n19023 = n19022 ^ n18934 ;
  assign n19024 = n19023 ^ n18938 ;
  assign n19025 = n19024 ^ n18934 ;
  assign n19026 = n19020 & ~n19025 ;
  assign n19027 = n19026 ^ n19023 ;
  assign n18936 = n18725 ^ n18724 ;
  assign n19199 = n19027 ^ n18936 ;
  assign n19200 = n19199 ^ n18631 ;
  assign n19201 = n18646 & ~n19200 ;
  assign n19202 = n19201 ^ n18631 ;
  assign n19204 = n19202 ^ n17791 ;
  assign n19203 = n19202 ^ n19193 ;
  assign n19205 = n19204 ^ n19203 ;
  assign n19206 = n19198 & ~n19205 ;
  assign n19207 = n19206 ^ n19204 ;
  assign n19416 = n19207 ^ n17825 ;
  assign n19417 = n19416 ^ x95 ;
  assign n19418 = n19417 ^ n19281 ;
  assign n19419 = n19418 ^ n19416 ;
  assign n19420 = ~n19415 & n19419 ;
  assign n19421 = n19420 ^ n19417 ;
  assign n19501 = n19421 ^ x94 ;
  assign n19500 = ~n19497 & n19499 ;
  assign n19533 = n19501 ^ n19500 ;
  assign n19543 = n19542 ^ n19533 ;
  assign n19630 = ~n18853 & n19543 ;
  assign n19534 = n18859 ^ n18854 ;
  assign n19631 = n19630 ^ n19534 ;
  assign n19711 = n19710 ^ n19631 ;
  assign n19712 = n19711 ^ x230 ;
  assign n19713 = n19712 ^ n19706 ;
  assign n19714 = n19713 ^ n19711 ;
  assign n19715 = n19709 & ~n19714 ;
  assign n19716 = n19715 ^ n19712 ;
  assign n19886 = n19716 ^ x229 ;
  assign n19887 = n19885 & ~n19886 ;
  assign n19632 = n19631 ^ n18217 ;
  assign n19642 = n19641 ^ n19631 ;
  assign n19643 = n19632 & ~n19642 ;
  assign n19644 = n19643 ^ n18217 ;
  assign n19717 = n19644 ^ n18212 ;
  assign n19535 = n19534 ^ n19533 ;
  assign n19544 = ~n19535 & ~n19543 ;
  assign n19545 = n19544 ^ n19534 ;
  assign n18937 = n18936 ^ n18934 ;
  assign n19028 = ~n18937 & n19027 ;
  assign n18935 = n18934 ^ n18652 ;
  assign n19029 = n19028 ^ n18935 ;
  assign n18933 = n18727 ^ n18726 ;
  assign n19030 = n19029 ^ n18933 ;
  assign n19031 = n19030 ^ n18652 ;
  assign n19032 = ~n17949 & n19031 ;
  assign n19033 = n19032 ^ n18652 ;
  assign n19209 = n19033 ^ n17825 ;
  assign n19208 = n19202 ^ n19033 ;
  assign n19210 = n19209 ^ n19208 ;
  assign n19211 = n19207 & ~n19210 ;
  assign n19212 = n19211 ^ n19209 ;
  assign n19422 = n19212 ^ n17320 ;
  assign n19424 = n19422 ^ x94 ;
  assign n19423 = n19422 ^ n19416 ;
  assign n19425 = n19424 ^ n19423 ;
  assign n19426 = ~n19421 & n19425 ;
  assign n19427 = n19426 ^ n19424 ;
  assign n19503 = n19427 ^ x93 ;
  assign n19502 = n19500 & n19501 ;
  assign n19529 = n19503 ^ n19502 ;
  assign n19546 = n19545 ^ n19529 ;
  assign n19627 = n18850 & n19546 ;
  assign n19530 = n18861 ^ n18850 ;
  assign n19531 = n19530 ^ n18849 ;
  assign n19628 = n19627 ^ n19531 ;
  assign n19718 = n19717 ^ n19628 ;
  assign n19720 = n19718 ^ x229 ;
  assign n19719 = n19718 ^ n19711 ;
  assign n19721 = n19720 ^ n19719 ;
  assign n19722 = n19716 & ~n19721 ;
  assign n19723 = n19722 ^ n19720 ;
  assign n19888 = n19723 ^ x228 ;
  assign n19889 = ~n19887 & n19888 ;
  assign n19629 = n19628 ^ n18212 ;
  assign n19645 = n19644 ^ n19628 ;
  assign n19646 = n19629 & n19645 ;
  assign n19647 = n19646 ^ n18212 ;
  assign n19724 = n19647 ^ n18209 ;
  assign n19532 = n19531 ^ n19529 ;
  assign n19547 = ~n19532 & ~n19546 ;
  assign n19548 = n19547 ^ n19531 ;
  assign n19034 = n19033 ^ n17320 ;
  assign n19213 = ~n19034 & ~n19212 ;
  assign n19214 = n19213 ^ n17320 ;
  assign n19428 = n19214 ^ n17341 ;
  assign n19220 = n18729 ^ n18728 ;
  assign n19215 = n18673 ^ n18652 ;
  assign n19216 = n19215 ^ n18673 ;
  assign n19217 = n19216 ^ n18933 ;
  assign n19218 = ~n19029 & ~n19217 ;
  assign n19219 = n19218 ^ n19215 ;
  assign n19221 = n19220 ^ n19219 ;
  assign n19222 = n19221 ^ n18673 ;
  assign n19223 = n17957 & n19222 ;
  assign n19224 = n19223 ^ n18673 ;
  assign n19429 = n19428 ^ n19224 ;
  assign n19431 = n19429 ^ x93 ;
  assign n19430 = n19429 ^ n19422 ;
  assign n19432 = n19431 ^ n19430 ;
  assign n19433 = ~n19427 & n19432 ;
  assign n19434 = n19433 ^ n19431 ;
  assign n19505 = n19434 ^ x92 ;
  assign n19504 = ~n19502 & ~n19503 ;
  assign n19526 = n19505 ^ n19504 ;
  assign n19549 = n19548 ^ n19526 ;
  assign n19624 = n18782 & n19549 ;
  assign n19527 = n18865 ^ n18846 ;
  assign n19625 = n19624 ^ n19527 ;
  assign n19725 = n19724 ^ n19625 ;
  assign n19727 = n19725 ^ x228 ;
  assign n19726 = n19725 ^ n19718 ;
  assign n19728 = n19727 ^ n19726 ;
  assign n19729 = n19723 & ~n19728 ;
  assign n19730 = n19729 ^ n19727 ;
  assign n19890 = n19730 ^ x227 ;
  assign n19891 = n19889 & ~n19890 ;
  assign n19626 = n19625 ^ n18209 ;
  assign n19648 = n19647 ^ n19625 ;
  assign n19649 = n19626 & ~n19648 ;
  assign n19650 = n19649 ^ n18209 ;
  assign n19731 = n19650 ^ n18204 ;
  assign n19528 = n19527 ^ n19526 ;
  assign n19550 = n19528 & ~n19549 ;
  assign n19551 = n19550 ^ n19527 ;
  assign n19225 = n19224 ^ n19214 ;
  assign n19226 = n19224 ^ n17341 ;
  assign n19227 = ~n19225 & n19226 ;
  assign n19228 = n19227 ^ n17341 ;
  assign n19435 = n19228 ^ n17480 ;
  assign n19230 = n19220 ^ n18673 ;
  assign n19231 = ~n19219 & ~n19230 ;
  assign n19232 = n19231 ^ n18673 ;
  assign n19229 = n18731 ^ n18730 ;
  assign n19233 = n19232 ^ n19229 ;
  assign n19234 = n17843 & ~n19233 ;
  assign n19235 = n19234 ^ n18756 ;
  assign n19436 = n19435 ^ n19235 ;
  assign n19438 = n19436 ^ x92 ;
  assign n19437 = n19436 ^ n19429 ;
  assign n19439 = n19438 ^ n19437 ;
  assign n19440 = ~n19434 & n19439 ;
  assign n19441 = n19440 ^ n19438 ;
  assign n19507 = n19441 ^ x91 ;
  assign n19506 = n19504 & ~n19505 ;
  assign n19522 = n19507 ^ n19506 ;
  assign n19552 = n19551 ^ n19522 ;
  assign n19621 = ~n18868 & ~n19552 ;
  assign n19523 = n18868 ^ n18686 ;
  assign n19524 = n19523 ^ n18867 ;
  assign n19622 = n19621 ^ n19524 ;
  assign n19732 = n19731 ^ n19622 ;
  assign n19734 = n19732 ^ x227 ;
  assign n19733 = n19732 ^ n19725 ;
  assign n19735 = n19734 ^ n19733 ;
  assign n19736 = ~n19730 & n19735 ;
  assign n19737 = n19736 ^ n19734 ;
  assign n19892 = n19737 ^ x226 ;
  assign n19893 = ~n19891 & ~n19892 ;
  assign n19623 = n19622 ^ n18204 ;
  assign n19651 = n19650 ^ n19622 ;
  assign n19652 = ~n19623 & ~n19651 ;
  assign n19653 = n19652 ^ n18204 ;
  assign n19738 = n19653 ^ n18200 ;
  assign n19525 = n19524 ^ n19522 ;
  assign n19553 = ~n19525 & n19552 ;
  assign n19554 = n19553 ^ n19524 ;
  assign n19236 = n19235 ^ n19228 ;
  assign n19237 = n19235 ^ n17480 ;
  assign n19238 = n19236 & ~n19237 ;
  assign n19239 = n19238 ^ n17480 ;
  assign n19442 = n19239 ^ n17572 ;
  assign n19246 = n18734 ^ n18732 ;
  assign n19240 = n18793 ^ n17974 ;
  assign n19241 = n19240 ^ n18756 ;
  assign n19242 = n19241 ^ n19229 ;
  assign n19243 = n19242 ^ n19240 ;
  assign n19244 = n19233 & n19243 ;
  assign n19245 = n19244 ^ n19241 ;
  assign n19247 = n19246 ^ n19245 ;
  assign n19248 = n19247 ^ n18793 ;
  assign n19249 = n17974 & ~n19248 ;
  assign n19250 = n19249 ^ n19247 ;
  assign n19443 = n19442 ^ n19250 ;
  assign n19445 = n19443 ^ x91 ;
  assign n19444 = n19443 ^ n19436 ;
  assign n19446 = n19445 ^ n19444 ;
  assign n19447 = n19441 & ~n19446 ;
  assign n19448 = n19447 ^ n19445 ;
  assign n19509 = n19448 ^ x90 ;
  assign n19508 = n19506 & n19507 ;
  assign n19520 = n19509 ^ n19508 ;
  assign n19555 = n19554 ^ n19520 ;
  assign n19618 = n18870 & n19555 ;
  assign n19619 = n19618 ^ n19063 ;
  assign n19739 = n19738 ^ n19619 ;
  assign n19741 = n19739 ^ x226 ;
  assign n19740 = n19739 ^ n19732 ;
  assign n19742 = n19741 ^ n19740 ;
  assign n19743 = n19737 & ~n19742 ;
  assign n19744 = n19743 ^ n19741 ;
  assign n19894 = n19744 ^ x225 ;
  assign n19895 = ~n19893 & ~n19894 ;
  assign n19620 = n19619 ^ n18200 ;
  assign n19654 = n19653 ^ n19619 ;
  assign n19655 = ~n19620 & n19654 ;
  assign n19656 = n19655 ^ n18200 ;
  assign n19745 = n19656 ^ n18196 ;
  assign n19521 = n19520 ^ n19063 ;
  assign n19556 = n19521 & ~n19555 ;
  assign n19557 = n19556 ^ n19063 ;
  assign n19251 = n19250 ^ n19239 ;
  assign n19252 = n19250 ^ n17572 ;
  assign n19253 = n19251 & n19252 ;
  assign n19254 = n19253 ^ n17572 ;
  assign n19449 = n19254 ^ n17684 ;
  assign n19257 = n19246 ^ n19240 ;
  assign n19258 = n19245 & n19257 ;
  assign n19256 = n19240 ^ n18813 ;
  assign n19259 = n19258 ^ n19256 ;
  assign n19255 = n18736 ^ n18735 ;
  assign n19260 = n19259 ^ n19255 ;
  assign n19261 = n19260 ^ n18813 ;
  assign n19262 = n17988 & ~n19261 ;
  assign n19263 = n19262 ^ n18813 ;
  assign n19450 = n19449 ^ n19263 ;
  assign n19452 = n19450 ^ x90 ;
  assign n19451 = n19450 ^ n19443 ;
  assign n19453 = n19452 ^ n19451 ;
  assign n19454 = ~n19448 & n19453 ;
  assign n19455 = n19454 ^ n19452 ;
  assign n19517 = n19455 ^ x89 ;
  assign n19510 = n19508 & ~n19509 ;
  assign n19518 = n19517 ^ n19510 ;
  assign n19558 = n19557 ^ n19518 ;
  assign n19657 = ~n18877 & n19558 ;
  assign n19658 = n19657 ^ n19070 ;
  assign n19746 = n19745 ^ n19658 ;
  assign n19748 = n19746 ^ x225 ;
  assign n19747 = n19746 ^ n19739 ;
  assign n19749 = n19748 ^ n19747 ;
  assign n19750 = ~n19744 & n19749 ;
  assign n19751 = n19750 ^ n19748 ;
  assign n19896 = n19751 ^ x224 ;
  assign n19897 = n19895 & ~n19896 ;
  assign n19659 = n19658 ^ n19656 ;
  assign n19660 = n19658 ^ n18196 ;
  assign n19661 = n19659 & ~n19660 ;
  assign n19662 = n19661 ^ n18196 ;
  assign n19752 = n19662 ^ n18246 ;
  assign n19519 = n19518 ^ n19070 ;
  assign n19559 = n19519 & ~n19558 ;
  assign n19560 = n19559 ^ n19070 ;
  assign n19513 = n19510 ^ n19450 ;
  assign n19514 = ~n19455 & n19513 ;
  assign n19511 = n19510 ^ n19455 ;
  assign n19512 = x89 & n19511 ;
  assign n19515 = n19514 ^ n19512 ;
  assign n19275 = n19255 ^ n18813 ;
  assign n19276 = n19259 & n19275 ;
  assign n19272 = n18738 ^ n18737 ;
  assign n19273 = n19272 ^ n19255 ;
  assign n19271 = n18843 ^ n18004 ;
  assign n19274 = n19273 ^ n19271 ;
  assign n19277 = n19276 ^ n19274 ;
  assign n19278 = n19277 ^ n18843 ;
  assign n19279 = n18004 & ~n19278 ;
  assign n19268 = n18843 ^ n17746 ;
  assign n19267 = n17684 ^ x88 ;
  assign n19269 = n19268 ^ n19267 ;
  assign n19264 = n19263 ^ n19254 ;
  assign n19265 = n19263 ^ n17684 ;
  assign n19266 = n19264 & ~n19265 ;
  assign n19270 = n19269 ^ n19266 ;
  assign n19280 = n19279 ^ n19270 ;
  assign n19516 = n19515 ^ n19280 ;
  assign n19561 = n19560 ^ n19516 ;
  assign n19615 = ~n18777 & n19561 ;
  assign n19616 = n19615 ^ n19079 ;
  assign n19753 = n19752 ^ n19616 ;
  assign n19755 = n19753 ^ x224 ;
  assign n19754 = n19753 ^ n19746 ;
  assign n19756 = n19755 ^ n19754 ;
  assign n19757 = ~n19751 & n19756 ;
  assign n19758 = n19757 ^ n19755 ;
  assign n19898 = n19758 ^ x239 ;
  assign n19899 = ~n19897 & n19898 ;
  assign n19617 = n19616 ^ n18246 ;
  assign n19663 = n19662 ^ n19616 ;
  assign n19664 = ~n19617 & ~n19663 ;
  assign n19665 = n19664 ^ n18246 ;
  assign n19759 = n19665 ^ n18191 ;
  assign n19567 = n18910 ^ x71 ;
  assign n19562 = n19087 ^ n19079 ;
  assign n19563 = n19562 ^ n19087 ;
  assign n19564 = n19563 ^ n19516 ;
  assign n19565 = ~n19561 & ~n19564 ;
  assign n19566 = n19565 ^ n19562 ;
  assign n19611 = n19567 ^ n19566 ;
  assign n19612 = n19611 ^ n19087 ;
  assign n19613 = n18774 & n19612 ;
  assign n19614 = n19613 ^ n19087 ;
  assign n19760 = n19759 ^ n19614 ;
  assign n19762 = n19760 ^ x239 ;
  assign n19761 = n19760 ^ n19753 ;
  assign n19763 = n19762 ^ n19761 ;
  assign n19764 = ~n19758 & n19763 ;
  assign n19765 = n19764 ^ n19762 ;
  assign n19900 = n19765 ^ x238 ;
  assign n19901 = ~n19899 & ~n19900 ;
  assign n19666 = n19665 ^ n19614 ;
  assign n18928 = n18896 ^ n18892 ;
  assign n19569 = n19087 ^ n18928 ;
  assign n19568 = n19567 ^ n18928 ;
  assign n19570 = n19569 ^ n19568 ;
  assign n19571 = n19566 & n19570 ;
  assign n19572 = n19571 ^ n19569 ;
  assign n18930 = n18911 ^ x70 ;
  assign n18931 = n18930 ^ n18909 ;
  assign n19606 = n19572 ^ n18931 ;
  assign n19607 = n19606 ^ n18892 ;
  assign n19608 = ~n18896 & n19607 ;
  assign n19609 = n19608 ^ n19606 ;
  assign n19667 = n19609 ^ n18191 ;
  assign n19668 = n19667 ^ n19614 ;
  assign n19669 = n19668 ^ n19609 ;
  assign n19670 = n19666 & n19669 ;
  assign n19671 = n19670 ^ n19667 ;
  assign n19766 = n19671 ^ n18187 ;
  assign n19768 = n19766 ^ x238 ;
  assign n19767 = n19766 ^ n19760 ;
  assign n19769 = n19768 ^ n19767 ;
  assign n19770 = ~n19765 & n19769 ;
  assign n19771 = n19770 ^ n19768 ;
  assign n19902 = n19771 ^ x237 ;
  assign n19903 = ~n19901 & ~n19902 ;
  assign n19610 = n19609 ^ n18187 ;
  assign n19672 = n19610 & n19671 ;
  assign n19673 = n19672 ^ n18187 ;
  assign n19772 = n19673 ^ n18258 ;
  assign n18932 = n18931 ^ n18928 ;
  assign n19573 = ~n18932 & ~n19572 ;
  assign n18929 = n18928 ^ n18902 ;
  assign n19574 = n19573 ^ n18929 ;
  assign n18926 = n18925 ^ x69 ;
  assign n19601 = n19574 ^ n18926 ;
  assign n19602 = n19601 ^ n18902 ;
  assign n19603 = n18894 & n19602 ;
  assign n19604 = n19603 ^ n18902 ;
  assign n19773 = n19772 ^ n19604 ;
  assign n19775 = n19773 ^ x237 ;
  assign n19774 = n19773 ^ n19766 ;
  assign n19776 = n19775 ^ n19774 ;
  assign n19777 = n19771 & ~n19776 ;
  assign n19778 = n19777 ^ n19775 ;
  assign n19904 = n19778 ^ x236 ;
  assign n19905 = n19903 & n19904 ;
  assign n19605 = n19604 ^ n18258 ;
  assign n19674 = n19673 ^ n19604 ;
  assign n19675 = n19605 & n19674 ;
  assign n19676 = n19675 ^ n18258 ;
  assign n19703 = n19676 ^ n18182 ;
  assign n18927 = n18926 ^ n18902 ;
  assign n19575 = ~n18927 & n19574 ;
  assign n19576 = n19575 ^ n18926 ;
  assign n19677 = n19576 ^ n19457 ;
  assign n19678 = n18955 & ~n19677 ;
  assign n19679 = n19678 ^ n18951 ;
  assign n19704 = n19703 ^ n19679 ;
  assign n19780 = n19704 ^ x236 ;
  assign n19779 = n19773 ^ n19704 ;
  assign n19781 = n19780 ^ n19779 ;
  assign n19782 = ~n19778 & n19781 ;
  assign n19783 = n19782 ^ n19780 ;
  assign n19906 = n19783 ^ x235 ;
  assign n19907 = n19905 & n19906 ;
  assign n19705 = n19704 ^ x235 ;
  assign n19784 = n19705 & ~n19783 ;
  assign n19785 = n19784 ^ x235 ;
  assign n19908 = n19785 ^ x234 ;
  assign n19680 = n19679 ^ n19676 ;
  assign n19681 = n19679 ^ n18182 ;
  assign n19682 = ~n19680 & ~n19681 ;
  assign n19683 = n19682 ^ n18182 ;
  assign n19786 = n19683 ^ n18266 ;
  assign n19584 = n19458 ^ n19457 ;
  assign n19577 = n18955 ^ n18951 ;
  assign n19578 = n19577 ^ n19576 ;
  assign n19579 = n19457 ^ n19114 ;
  assign n19580 = n19579 ^ n19114 ;
  assign n19581 = n19580 ^ n19576 ;
  assign n19582 = n19578 & n19581 ;
  assign n19583 = n19582 ^ n19579 ;
  assign n19596 = n19584 ^ n19583 ;
  assign n19597 = n19596 ^ n19114 ;
  assign n19598 = ~n18953 & ~n19597 ;
  assign n19599 = n19598 ^ n19114 ;
  assign n19787 = n19786 ^ n19599 ;
  assign n19909 = n19908 ^ n19787 ;
  assign n19910 = n19907 & n19909 ;
  assign n19788 = n19787 ^ n19785 ;
  assign n19600 = n19599 ^ n18266 ;
  assign n19684 = n19683 ^ n19599 ;
  assign n19685 = n19600 & ~n19684 ;
  assign n19686 = n19685 ^ n18266 ;
  assign n19789 = n19686 ^ n18177 ;
  assign n19590 = n19460 ^ n19459 ;
  assign n19586 = n19122 ^ n19114 ;
  assign n19585 = n19584 ^ n19122 ;
  assign n19587 = n19586 ^ n19585 ;
  assign n19588 = n19583 & ~n19587 ;
  assign n19589 = n19588 ^ n19586 ;
  assign n19591 = n19590 ^ n19589 ;
  assign n19592 = n19591 ^ n19122 ;
  assign n19593 = ~n18770 & n19592 ;
  assign n19594 = n19593 ^ n19122 ;
  assign n19790 = n19789 ^ n19594 ;
  assign n19791 = n19790 ^ x234 ;
  assign n19792 = n19791 ^ n19785 ;
  assign n19793 = n19792 ^ n19790 ;
  assign n19794 = ~n19788 & n19793 ;
  assign n19795 = n19794 ^ n19791 ;
  assign n19911 = n19795 ^ x233 ;
  assign n19912 = n19910 & ~n19911 ;
  assign n19696 = n19462 ^ n19461 ;
  assign n19692 = n19130 ^ n19122 ;
  assign n19691 = n19590 ^ n19130 ;
  assign n19693 = n19692 ^ n19691 ;
  assign n19694 = n19589 & n19693 ;
  assign n19695 = n19694 ^ n19692 ;
  assign n19697 = n19696 ^ n19695 ;
  assign n19698 = n19697 ^ n19130 ;
  assign n19699 = ~n18970 & n19698 ;
  assign n19700 = n19699 ^ n19130 ;
  assign n19595 = n19594 ^ n18177 ;
  assign n19687 = n19686 ^ n19594 ;
  assign n19688 = ~n19595 & ~n19687 ;
  assign n19689 = n19688 ^ n18177 ;
  assign n19690 = n19689 ^ n17879 ;
  assign n19701 = n19700 ^ n19690 ;
  assign n19797 = n19701 ^ x233 ;
  assign n19796 = n19790 ^ n19701 ;
  assign n19798 = n19797 ^ n19796 ;
  assign n19799 = n19795 & ~n19798 ;
  assign n19800 = n19799 ^ n19797 ;
  assign n19913 = n19800 ^ x232 ;
  assign n19914 = n19912 & n19913 ;
  assign n19702 = n19701 ^ x232 ;
  assign n19801 = n19702 & ~n19800 ;
  assign n19802 = n19801 ^ x232 ;
  assign n19915 = n19802 ^ x247 ;
  assign n19803 = n19700 ^ n19689 ;
  assign n19810 = n19463 ^ n19456 ;
  assign n19804 = n18980 ^ n18976 ;
  assign n19806 = n19804 ^ n19130 ;
  assign n19805 = n19804 ^ n19696 ;
  assign n19807 = n19806 ^ n19805 ;
  assign n19808 = ~n19695 & ~n19807 ;
  assign n19809 = n19808 ^ n19806 ;
  assign n19811 = n19810 ^ n19809 ;
  assign n19812 = n19811 ^ n19804 ;
  assign n19813 = n18979 & ~n19812 ;
  assign n19814 = n19813 ^ n19804 ;
  assign n19815 = n19814 ^ n17879 ;
  assign n19816 = n19815 ^ n19689 ;
  assign n19817 = n19816 ^ n19814 ;
  assign n19818 = ~n19803 & ~n19817 ;
  assign n19819 = n19818 ^ n19815 ;
  assign n19820 = n19819 ^ n17858 ;
  assign n19916 = n19915 ^ n19820 ;
  assign n19917 = ~n19914 & n19916 ;
  assign n19821 = n19820 ^ n19802 ;
  assign n19830 = n19814 ^ n17858 ;
  assign n19831 = n19819 & ~n19830 ;
  assign n19832 = n19831 ^ n17858 ;
  assign n19833 = n19832 ^ n18173 ;
  assign n19822 = n19465 ^ n19464 ;
  assign n19824 = n19822 ^ n19804 ;
  assign n19823 = n19822 ^ n19810 ;
  assign n19825 = n19824 ^ n19823 ;
  assign n19826 = n19809 & ~n19825 ;
  assign n19827 = n19826 ^ n19824 ;
  assign n19828 = ~n18985 & ~n19827 ;
  assign n19829 = n19828 ^ n18984 ;
  assign n19834 = n19833 ^ n19829 ;
  assign n19835 = n19834 ^ x247 ;
  assign n19836 = n19835 ^ n19802 ;
  assign n19837 = n19836 ^ n19834 ;
  assign n19838 = n19821 & n19837 ;
  assign n19839 = n19838 ^ n19835 ;
  assign n19918 = n19839 ^ x246 ;
  assign n19919 = n19917 & ~n19918 ;
  assign n19850 = n19832 ^ n19829 ;
  assign n19851 = n19833 & ~n19850 ;
  assign n19852 = n19851 ^ n18173 ;
  assign n19853 = n19852 ^ n17897 ;
  assign n19845 = n19467 ^ n19466 ;
  assign n19843 = n19822 ^ n19148 ;
  assign n19840 = n18985 ^ n18984 ;
  assign n19841 = n19840 ^ n19822 ;
  assign n19842 = n19827 & n19841 ;
  assign n19844 = n19843 ^ n19842 ;
  assign n19846 = n19845 ^ n19844 ;
  assign n19847 = n19846 ^ n19148 ;
  assign n19848 = ~n18988 & n19847 ;
  assign n19849 = n19848 ^ n19148 ;
  assign n19854 = n19853 ^ n19849 ;
  assign n19856 = n19854 ^ x246 ;
  assign n19855 = n19854 ^ n19834 ;
  assign n19857 = n19856 ^ n19855 ;
  assign n19858 = ~n19839 & n19857 ;
  assign n19859 = n19858 ^ n19856 ;
  assign n19881 = n19859 ^ x245 ;
  assign n19922 = n19919 ^ n19881 ;
  assign n20463 = n19923 ^ n19922 ;
  assign n19929 = n18741 & ~n19922 ;
  assign n19930 = n19929 ^ n19536 ;
  assign n19934 = n19930 ^ n17727 ;
  assign n19935 = x391 & n19934 ;
  assign n20396 = n19935 ^ x390 ;
  assign n19931 = n17727 & n19930 ;
  assign n19932 = n19931 ^ n18742 ;
  assign n19927 = n19539 ^ n19538 ;
  assign n19924 = n19922 & n19923 ;
  assign n19920 = ~n19881 & n19919 ;
  assign n19869 = n19469 ^ n19468 ;
  assign n19865 = n19156 ^ n19148 ;
  assign n19864 = n19845 ^ n19156 ;
  assign n19866 = n19865 ^ n19864 ;
  assign n19867 = ~n19844 & ~n19866 ;
  assign n19868 = n19867 ^ n19865 ;
  assign n19870 = n19869 ^ n19868 ;
  assign n19871 = n19870 ^ n19156 ;
  assign n19872 = n18991 & ~n19871 ;
  assign n19873 = n19872 ^ n19156 ;
  assign n19860 = n19852 ^ n19849 ;
  assign n19861 = n19853 & ~n19860 ;
  assign n19862 = n19861 ^ n17897 ;
  assign n19863 = n19862 ^ n17788 ;
  assign n19874 = n19873 ^ n19863 ;
  assign n19876 = n19874 ^ x245 ;
  assign n19875 = n19874 ^ n19854 ;
  assign n19877 = n19876 ^ n19875 ;
  assign n19878 = ~n19859 & n19877 ;
  assign n19879 = n19878 ^ n19876 ;
  assign n19880 = n19879 ^ x244 ;
  assign n19921 = n19920 ^ n19880 ;
  assign n19925 = n19924 ^ n19921 ;
  assign n19926 = n18769 & n19925 ;
  assign n19928 = n19927 ^ n19926 ;
  assign n19933 = n19932 ^ n19928 ;
  assign n20397 = n20396 ^ n19933 ;
  assign n19936 = n19935 ^ n19933 ;
  assign n19969 = n19931 ^ n19928 ;
  assign n19970 = n19932 & n19969 ;
  assign n19971 = n19970 ^ n18742 ;
  assign n19972 = n19971 ^ n18853 ;
  assign n19966 = n19542 ^ n19534 ;
  assign n19967 = n19966 ^ n19533 ;
  assign n19962 = ~n19880 & n19920 ;
  assign n19950 = n19471 ^ n19470 ;
  assign n19946 = n19164 ^ n19156 ;
  assign n19945 = n19869 ^ n19164 ;
  assign n19947 = n19946 ^ n19945 ;
  assign n19948 = n19868 & ~n19947 ;
  assign n19949 = n19948 ^ n19946 ;
  assign n19951 = n19950 ^ n19949 ;
  assign n19952 = n19951 ^ n19164 ;
  assign n19953 = n18942 & n19952 ;
  assign n19954 = n19953 ^ n19164 ;
  assign n19940 = n19873 ^ n17788 ;
  assign n19941 = n19873 ^ n19862 ;
  assign n19942 = n19940 & ~n19941 ;
  assign n19943 = n19942 ^ n17788 ;
  assign n19944 = n19943 ^ n17911 ;
  assign n19955 = n19954 ^ n19944 ;
  assign n19957 = n19955 ^ x244 ;
  assign n19956 = n19955 ^ n19874 ;
  assign n19958 = n19957 ^ n19956 ;
  assign n19959 = ~n19879 & n19958 ;
  assign n19960 = n19959 ^ n19957 ;
  assign n19961 = n19960 ^ x243 ;
  assign n19963 = n19962 ^ n19961 ;
  assign n19937 = n19927 ^ n19924 ;
  assign n19938 = ~n19925 & ~n19937 ;
  assign n19939 = n19938 ^ n19927 ;
  assign n19964 = n19963 ^ n19939 ;
  assign n19965 = ~n19534 & ~n19964 ;
  assign n19968 = n19967 ^ n19965 ;
  assign n19973 = n19972 ^ n19968 ;
  assign n19974 = n19973 ^ x390 ;
  assign n19975 = n19974 ^ n19933 ;
  assign n19976 = n19975 ^ n19973 ;
  assign n19977 = n19936 & ~n19976 ;
  assign n19978 = n19977 ^ n19974 ;
  assign n20398 = n19978 ^ x389 ;
  assign n20399 = ~n20397 & n20398 ;
  assign n20012 = n19971 ^ n19968 ;
  assign n20013 = ~n19972 & n20012 ;
  assign n20014 = n20013 ^ n18853 ;
  assign n20015 = n20014 ^ n18850 ;
  assign n20009 = n19545 ^ n19531 ;
  assign n20010 = n20009 ^ n19529 ;
  assign n20005 = ~n19961 & ~n19962 ;
  assign n19993 = n19473 ^ n19472 ;
  assign n19989 = n19172 ^ n19164 ;
  assign n19988 = n19950 ^ n19172 ;
  assign n19990 = n19989 ^ n19988 ;
  assign n19991 = n19949 & n19990 ;
  assign n19992 = n19991 ^ n19989 ;
  assign n19994 = n19993 ^ n19992 ;
  assign n19995 = n19994 ^ n19172 ;
  assign n19996 = n18300 & ~n19995 ;
  assign n19997 = n19996 ^ n19172 ;
  assign n19983 = n19954 ^ n17911 ;
  assign n19984 = n19954 ^ n19943 ;
  assign n19985 = ~n19983 & ~n19984 ;
  assign n19986 = n19985 ^ n17911 ;
  assign n19987 = n19986 ^ n17853 ;
  assign n19998 = n19997 ^ n19987 ;
  assign n20000 = n19998 ^ x243 ;
  assign n19999 = n19998 ^ n19955 ;
  assign n20001 = n20000 ^ n19999 ;
  assign n20002 = n19960 & ~n20001 ;
  assign n20003 = n20002 ^ n20000 ;
  assign n20004 = n20003 ^ x242 ;
  assign n20006 = n20005 ^ n20004 ;
  assign n19979 = n19967 ^ n19963 ;
  assign n19980 = n19967 ^ n19939 ;
  assign n19981 = ~n19979 & ~n19980 ;
  assign n19982 = n19981 ^ n19963 ;
  assign n20007 = n20006 ^ n19982 ;
  assign n20008 = n19531 & ~n20007 ;
  assign n20011 = n20010 ^ n20008 ;
  assign n20016 = n20015 ^ n20011 ;
  assign n20018 = n20016 ^ x389 ;
  assign n20017 = n20016 ^ n19973 ;
  assign n20019 = n20018 ^ n20017 ;
  assign n20020 = ~n19978 & n20019 ;
  assign n20021 = n20020 ^ n20018 ;
  assign n20400 = n20021 ^ x388 ;
  assign n20401 = ~n20399 & n20400 ;
  assign n20053 = n20014 ^ n20011 ;
  assign n20054 = ~n20015 & n20053 ;
  assign n20055 = n20054 ^ n18850 ;
  assign n20056 = n20055 ^ n18782 ;
  assign n20050 = n19548 ^ n19527 ;
  assign n20051 = n20050 ^ n19526 ;
  assign n20046 = ~n20004 & ~n20005 ;
  assign n20042 = n19998 ^ x242 ;
  assign n20043 = ~n20003 & n20042 ;
  assign n20044 = n20043 ^ x242 ;
  assign n20035 = n19475 ^ n19474 ;
  assign n20031 = n19180 ^ n19172 ;
  assign n20030 = n19993 ^ n19180 ;
  assign n20032 = n20031 ^ n20030 ;
  assign n20033 = n19992 & ~n20032 ;
  assign n20034 = n20033 ^ n20031 ;
  assign n20036 = n20035 ^ n20034 ;
  assign n20037 = n20036 ^ n19180 ;
  assign n20038 = ~n18448 & ~n20037 ;
  assign n20039 = n20038 ^ n19180 ;
  assign n20025 = n19997 ^ n17853 ;
  assign n20026 = n19997 ^ n19986 ;
  assign n20027 = ~n20025 & n20026 ;
  assign n20028 = n20027 ^ n17853 ;
  assign n20029 = n20028 ^ n17923 ;
  assign n20040 = n20039 ^ n20029 ;
  assign n20041 = n20040 ^ x241 ;
  assign n20045 = n20044 ^ n20041 ;
  assign n20047 = n20046 ^ n20045 ;
  assign n20022 = n20010 ^ n20006 ;
  assign n20023 = n20007 & ~n20022 ;
  assign n20024 = n20023 ^ n20010 ;
  assign n20048 = n20047 ^ n20024 ;
  assign n20049 = n19527 & ~n20048 ;
  assign n20052 = n20051 ^ n20049 ;
  assign n20057 = n20056 ^ n20052 ;
  assign n20059 = n20057 ^ x388 ;
  assign n20058 = n20057 ^ n20016 ;
  assign n20060 = n20059 ^ n20058 ;
  assign n20061 = n20021 & ~n20060 ;
  assign n20062 = n20061 ^ n20059 ;
  assign n20402 = n20062 ^ x387 ;
  assign n20403 = ~n20401 & n20402 ;
  assign n20096 = n20055 ^ n20052 ;
  assign n20097 = n20056 & ~n20096 ;
  assign n20098 = n20097 ^ n18782 ;
  assign n20099 = n20098 ^ n18868 ;
  assign n20093 = n19551 ^ n19524 ;
  assign n20094 = n20093 ^ n19522 ;
  assign n20089 = n20045 & n20046 ;
  assign n20066 = n20044 ^ n20040 ;
  assign n20078 = n20039 ^ n17923 ;
  assign n20079 = n20039 ^ n20028 ;
  assign n20080 = n20078 & ~n20079 ;
  assign n20081 = n20080 ^ n17923 ;
  assign n20072 = n19477 ^ n19476 ;
  assign n20068 = n19187 ^ n19180 ;
  assign n20067 = n20035 ^ n19187 ;
  assign n20069 = n20068 ^ n20067 ;
  assign n20070 = ~n20034 & n20069 ;
  assign n20071 = n20070 ^ n20068 ;
  assign n20073 = n20072 ^ n20071 ;
  assign n20074 = n20073 ^ n19187 ;
  assign n20075 = n18462 & ~n20074 ;
  assign n20076 = n20075 ^ n19187 ;
  assign n20077 = n20076 ^ n17931 ;
  assign n20082 = n20081 ^ n20077 ;
  assign n20083 = n20082 ^ x241 ;
  assign n20084 = n20083 ^ n20082 ;
  assign n20085 = n20084 ^ n20044 ;
  assign n20086 = n20066 & n20085 ;
  assign n20087 = n20086 ^ n20083 ;
  assign n20088 = n20087 ^ x240 ;
  assign n20090 = n20089 ^ n20088 ;
  assign n20063 = n20051 ^ n20047 ;
  assign n20064 = n20048 & ~n20063 ;
  assign n20065 = n20064 ^ n20051 ;
  assign n20091 = n20090 ^ n20065 ;
  assign n20092 = n19524 & ~n20091 ;
  assign n20095 = n20094 ^ n20092 ;
  assign n20100 = n20099 ^ n20095 ;
  assign n20102 = n20100 ^ x387 ;
  assign n20101 = n20100 ^ n20057 ;
  assign n20103 = n20102 ^ n20101 ;
  assign n20104 = ~n20062 & n20103 ;
  assign n20105 = n20104 ^ n20102 ;
  assign n20404 = n20105 ^ x386 ;
  assign n20405 = n20403 & n20404 ;
  assign n20140 = n20098 ^ n20095 ;
  assign n20141 = ~n20099 & n20140 ;
  assign n20142 = n20141 ^ n18868 ;
  assign n20143 = n20142 ^ n18870 ;
  assign n20137 = n19554 ^ n19063 ;
  assign n20138 = n20137 ^ n19520 ;
  assign n20133 = n20088 & ~n20089 ;
  assign n20114 = n20081 ^ n20076 ;
  assign n20121 = n19479 ^ n19478 ;
  assign n20115 = n19022 ^ n19020 ;
  assign n20117 = n20115 ^ n19187 ;
  assign n20116 = n20115 ^ n20072 ;
  assign n20118 = n20117 ^ n20116 ;
  assign n20119 = ~n20071 & n20118 ;
  assign n20120 = n20119 ^ n20117 ;
  assign n20122 = n20121 ^ n20120 ;
  assign n20123 = n20122 ^ n19020 ;
  assign n20124 = n19022 & n20123 ;
  assign n20125 = n20124 ^ n19020 ;
  assign n20126 = n20125 ^ n17931 ;
  assign n20127 = n20126 ^ n20076 ;
  assign n20128 = n20127 ^ n20125 ;
  assign n20129 = n20114 & ~n20128 ;
  assign n20130 = n20129 ^ n20126 ;
  assign n20131 = n20130 ^ n17848 ;
  assign n20110 = n20082 ^ x240 ;
  assign n20111 = ~n20087 & n20110 ;
  assign n20112 = n20111 ^ x240 ;
  assign n20113 = n20112 ^ x255 ;
  assign n20132 = n20131 ^ n20113 ;
  assign n20134 = n20133 ^ n20132 ;
  assign n20106 = n20094 ^ n20090 ;
  assign n20107 = n20094 ^ n20065 ;
  assign n20108 = n20106 & n20107 ;
  assign n20109 = n20108 ^ n20090 ;
  assign n20135 = n20134 ^ n20109 ;
  assign n20136 = n19063 & n20135 ;
  assign n20139 = n20138 ^ n20136 ;
  assign n20144 = n20143 ^ n20139 ;
  assign n20146 = n20144 ^ x386 ;
  assign n20145 = n20144 ^ n20100 ;
  assign n20147 = n20146 ^ n20145 ;
  assign n20148 = ~n20105 & n20147 ;
  assign n20149 = n20148 ^ n20146 ;
  assign n20406 = n20149 ^ x385 ;
  assign n20407 = n20405 & ~n20406 ;
  assign n20179 = n20142 ^ n20139 ;
  assign n20180 = ~n20143 & n20179 ;
  assign n20181 = n20180 ^ n18870 ;
  assign n20182 = n20181 ^ n18877 ;
  assign n20176 = n19557 ^ n19070 ;
  assign n20177 = n20176 ^ n19518 ;
  assign n20172 = ~n20132 & ~n20133 ;
  assign n20153 = n20131 ^ n20112 ;
  assign n20159 = n20121 ^ n20115 ;
  assign n20160 = ~n20120 & ~n20159 ;
  assign n20161 = n20160 ^ n20115 ;
  assign n20158 = n19482 ^ n19480 ;
  assign n20162 = n20161 ^ n20158 ;
  assign n20163 = n18934 & n20162 ;
  assign n20164 = n20163 ^ n19199 ;
  assign n20154 = n20125 ^ n17848 ;
  assign n20155 = ~n20130 & ~n20154 ;
  assign n20156 = n20155 ^ n17848 ;
  assign n20157 = n20156 ^ n18646 ;
  assign n20165 = n20164 ^ n20157 ;
  assign n20166 = n20165 ^ x255 ;
  assign n20167 = n20166 ^ n20112 ;
  assign n20168 = n20167 ^ n20165 ;
  assign n20169 = ~n20153 & n20168 ;
  assign n20170 = n20169 ^ n20166 ;
  assign n20171 = n20170 ^ x254 ;
  assign n20173 = n20172 ^ n20171 ;
  assign n20150 = n20138 ^ n20134 ;
  assign n20151 = ~n20135 & ~n20150 ;
  assign n20152 = n20151 ^ n20138 ;
  assign n20174 = n20173 ^ n20152 ;
  assign n20175 = n19070 & ~n20174 ;
  assign n20178 = n20177 ^ n20175 ;
  assign n20183 = n20182 ^ n20178 ;
  assign n20185 = n20183 ^ x385 ;
  assign n20184 = n20183 ^ n20144 ;
  assign n20186 = n20185 ^ n20184 ;
  assign n20187 = n20149 & ~n20186 ;
  assign n20188 = n20187 ^ n20185 ;
  assign n20408 = n20188 ^ x384 ;
  assign n20409 = ~n20407 & n20408 ;
  assign n20222 = n20181 ^ n20178 ;
  assign n20223 = ~n20182 & ~n20222 ;
  assign n20224 = n20223 ^ n18877 ;
  assign n20225 = n20224 ^ n18777 ;
  assign n20219 = n19560 ^ n19079 ;
  assign n20220 = n20219 ^ n19516 ;
  assign n20215 = n20171 & n20172 ;
  assign n20203 = n19484 ^ n19483 ;
  assign n20199 = n19199 ^ n19030 ;
  assign n20198 = n20161 ^ n19030 ;
  assign n20200 = n20199 ^ n20198 ;
  assign n20201 = ~n20162 & n20200 ;
  assign n20202 = n20201 ^ n20199 ;
  assign n20204 = n20203 ^ n20202 ;
  assign n20205 = n20204 ^ n19030 ;
  assign n20206 = ~n18652 & ~n20205 ;
  assign n20207 = n20206 ^ n19030 ;
  assign n20193 = n20164 ^ n20156 ;
  assign n20194 = n20164 ^ n18646 ;
  assign n20195 = n20193 & ~n20194 ;
  assign n20196 = n20195 ^ n18646 ;
  assign n20197 = n20196 ^ n17949 ;
  assign n20208 = n20207 ^ n20197 ;
  assign n20210 = n20208 ^ x254 ;
  assign n20209 = n20208 ^ n20165 ;
  assign n20211 = n20210 ^ n20209 ;
  assign n20212 = n20170 & ~n20211 ;
  assign n20213 = n20212 ^ n20210 ;
  assign n20214 = n20213 ^ x253 ;
  assign n20216 = n20215 ^ n20214 ;
  assign n20189 = n20177 ^ n20173 ;
  assign n20190 = n20177 ^ n20152 ;
  assign n20191 = ~n20189 & ~n20190 ;
  assign n20192 = n20191 ^ n20173 ;
  assign n20217 = n20216 ^ n20192 ;
  assign n20218 = ~n19079 & ~n20217 ;
  assign n20221 = n20220 ^ n20218 ;
  assign n20226 = n20225 ^ n20221 ;
  assign n20228 = n20226 ^ x384 ;
  assign n20227 = n20226 ^ n20183 ;
  assign n20229 = n20228 ^ n20227 ;
  assign n20230 = n20188 & ~n20229 ;
  assign n20231 = n20230 ^ n20228 ;
  assign n20410 = n20231 ^ x399 ;
  assign n20411 = ~n20409 & ~n20410 ;
  assign n20262 = n20224 ^ n20221 ;
  assign n20263 = n20225 & ~n20262 ;
  assign n20264 = n20263 ^ n18777 ;
  assign n20265 = n20264 ^ n18774 ;
  assign n20257 = ~n20214 & n20215 ;
  assign n20245 = n19486 ^ n19485 ;
  assign n20241 = n19221 ^ n19030 ;
  assign n20240 = n20203 ^ n19221 ;
  assign n20242 = n20241 ^ n20240 ;
  assign n20243 = n20202 & ~n20242 ;
  assign n20244 = n20243 ^ n20241 ;
  assign n20246 = n20245 ^ n20244 ;
  assign n20247 = n20246 ^ n19221 ;
  assign n20248 = n18673 & ~n20247 ;
  assign n20249 = n20248 ^ n19221 ;
  assign n20235 = n20207 ^ n20196 ;
  assign n20236 = n20207 ^ n17949 ;
  assign n20237 = n20235 & n20236 ;
  assign n20238 = n20237 ^ n17949 ;
  assign n20239 = n20238 ^ n17957 ;
  assign n20250 = n20249 ^ n20239 ;
  assign n20252 = n20250 ^ x253 ;
  assign n20251 = n20250 ^ n20208 ;
  assign n20253 = n20252 ^ n20251 ;
  assign n20254 = ~n20213 & n20253 ;
  assign n20255 = n20254 ^ n20252 ;
  assign n20256 = n20255 ^ x252 ;
  assign n20258 = n20257 ^ n20256 ;
  assign n20232 = n20220 ^ n20216 ;
  assign n20233 = n20217 & ~n20232 ;
  assign n20234 = n20233 ^ n20220 ;
  assign n20259 = n20258 ^ n20234 ;
  assign n20260 = ~n19087 & ~n20259 ;
  assign n20261 = n20260 ^ n19611 ;
  assign n20266 = n20265 ^ n20261 ;
  assign n20268 = n20266 ^ x399 ;
  assign n20267 = n20266 ^ n20226 ;
  assign n20269 = n20268 ^ n20267 ;
  assign n20270 = n20231 & ~n20269 ;
  assign n20271 = n20270 ^ n20268 ;
  assign n20412 = n20271 ^ x398 ;
  assign n20413 = n20411 & n20412 ;
  assign n20304 = n20264 ^ n20261 ;
  assign n20305 = ~n20265 & ~n20304 ;
  assign n20306 = n20305 ^ n18774 ;
  assign n20307 = n20306 ^ n18896 ;
  assign n20298 = n20258 ^ n19611 ;
  assign n20299 = n20259 & ~n20298 ;
  assign n20300 = n20299 ^ n19611 ;
  assign n20296 = ~n20256 & ~n20257 ;
  assign n20284 = n19488 ^ n19487 ;
  assign n20277 = n19229 ^ n18756 ;
  assign n20278 = n20277 ^ n19232 ;
  assign n20280 = n20278 ^ n19221 ;
  assign n20279 = n20278 ^ n20245 ;
  assign n20281 = n20280 ^ n20279 ;
  assign n20282 = ~n20244 & n20281 ;
  assign n20283 = n20282 ^ n20280 ;
  assign n20285 = n20284 ^ n20283 ;
  assign n20286 = n20285 ^ n20278 ;
  assign n20287 = ~n18756 & n20286 ;
  assign n20288 = n20287 ^ n20278 ;
  assign n20272 = n20249 ^ n20238 ;
  assign n20273 = n20249 ^ n17957 ;
  assign n20274 = n20272 & n20273 ;
  assign n20275 = n20274 ^ n17957 ;
  assign n20276 = n20275 ^ n17843 ;
  assign n20289 = n20288 ^ n20276 ;
  assign n20291 = n20289 ^ x252 ;
  assign n20290 = n20289 ^ n20250 ;
  assign n20292 = n20291 ^ n20290 ;
  assign n20293 = n20255 & ~n20292 ;
  assign n20294 = n20293 ^ n20291 ;
  assign n20295 = n20294 ^ x251 ;
  assign n20297 = n20296 ^ n20295 ;
  assign n20301 = n20300 ^ n20297 ;
  assign n20302 = n18928 & ~n20301 ;
  assign n20303 = n20302 ^ n19606 ;
  assign n20308 = n20307 ^ n20303 ;
  assign n20310 = n20308 ^ x398 ;
  assign n20309 = n20308 ^ n20266 ;
  assign n20311 = n20310 ^ n20309 ;
  assign n20312 = ~n20271 & n20311 ;
  assign n20313 = n20312 ^ n20310 ;
  assign n20414 = n20313 ^ x397 ;
  assign n20415 = ~n20413 & ~n20414 ;
  assign n20343 = n20306 ^ n20303 ;
  assign n20344 = n20307 & ~n20343 ;
  assign n20345 = n20344 ^ n18896 ;
  assign n20346 = n20345 ^ n18894 ;
  assign n20338 = n20295 & n20296 ;
  assign n20324 = n20284 ^ n20278 ;
  assign n20325 = n20283 & n20324 ;
  assign n20323 = n20278 ^ n19247 ;
  assign n20326 = n20325 ^ n20323 ;
  assign n20322 = n19490 ^ n19489 ;
  assign n20327 = n20326 ^ n20322 ;
  assign n20328 = n20327 ^ n19247 ;
  assign n20329 = ~n19240 & n20328 ;
  assign n20330 = n20329 ^ n19247 ;
  assign n20317 = n20288 ^ n20275 ;
  assign n20318 = n20288 ^ n17843 ;
  assign n20319 = ~n20317 & n20318 ;
  assign n20320 = n20319 ^ n17843 ;
  assign n20321 = n20320 ^ n17974 ;
  assign n20331 = n20330 ^ n20321 ;
  assign n20333 = n20331 ^ x251 ;
  assign n20332 = n20331 ^ n20289 ;
  assign n20334 = n20333 ^ n20332 ;
  assign n20335 = ~n20294 & n20334 ;
  assign n20336 = n20335 ^ n20333 ;
  assign n20337 = n20336 ^ x250 ;
  assign n20339 = n20338 ^ n20337 ;
  assign n20314 = n20300 ^ n19606 ;
  assign n20315 = n20301 & ~n20314 ;
  assign n20316 = n20315 ^ n19606 ;
  assign n20340 = n20339 ^ n20316 ;
  assign n20341 = ~n18902 & ~n20340 ;
  assign n20342 = n20341 ^ n19601 ;
  assign n20347 = n20346 ^ n20342 ;
  assign n20349 = n20347 ^ x397 ;
  assign n20348 = n20347 ^ n20308 ;
  assign n20350 = n20349 ^ n20348 ;
  assign n20351 = ~n20313 & n20350 ;
  assign n20352 = n20351 ^ n20349 ;
  assign n20416 = n20352 ^ x396 ;
  assign n20417 = n20415 & n20416 ;
  assign n20385 = n20345 ^ n20342 ;
  assign n20386 = n20346 & n20385 ;
  assign n20387 = n20386 ^ n18894 ;
  assign n20388 = n20387 ^ n18955 ;
  assign n20382 = n19577 ^ n19457 ;
  assign n20383 = n20382 ^ n19576 ;
  assign n20378 = ~n20337 & ~n20338 ;
  assign n20366 = n19492 ^ n19491 ;
  assign n20361 = n19260 ^ n19247 ;
  assign n20362 = n20361 ^ n19260 ;
  assign n20363 = n20362 ^ n20322 ;
  assign n20364 = ~n20326 & ~n20363 ;
  assign n20365 = n20364 ^ n20361 ;
  assign n20367 = n20366 ^ n20365 ;
  assign n20368 = n20367 ^ n19260 ;
  assign n20369 = n18813 & n20368 ;
  assign n20370 = n20369 ^ n19260 ;
  assign n20356 = n20330 ^ n20320 ;
  assign n20357 = n20330 ^ n17974 ;
  assign n20358 = n20356 & n20357 ;
  assign n20359 = n20358 ^ n17974 ;
  assign n20360 = n20359 ^ n17988 ;
  assign n20371 = n20370 ^ n20360 ;
  assign n20373 = n20371 ^ x250 ;
  assign n20372 = n20371 ^ n20331 ;
  assign n20374 = n20373 ^ n20372 ;
  assign n20375 = ~n20336 & n20374 ;
  assign n20376 = n20375 ^ n20373 ;
  assign n20377 = n20376 ^ x249 ;
  assign n20379 = n20378 ^ n20377 ;
  assign n20353 = n20339 ^ n19601 ;
  assign n20354 = n20340 & n20353 ;
  assign n20355 = n20354 ^ n19601 ;
  assign n20380 = n20379 ^ n20355 ;
  assign n20381 = ~n19577 & ~n20380 ;
  assign n20384 = n20383 ^ n20381 ;
  assign n20389 = n20388 ^ n20384 ;
  assign n20391 = n20389 ^ x396 ;
  assign n20390 = n20389 ^ n20347 ;
  assign n20392 = n20391 ^ n20390 ;
  assign n20393 = n20352 & ~n20392 ;
  assign n20394 = n20393 ^ n20391 ;
  assign n20395 = n20394 ^ x395 ;
  assign n20418 = n20417 ^ n20395 ;
  assign n20419 = n20418 ^ n19536 ;
  assign n20469 = x167 & n20419 ;
  assign n20464 = n20418 & n20463 ;
  assign n20461 = ~n20395 & ~n20417 ;
  assign n20450 = n20387 ^ n20384 ;
  assign n20451 = n20388 & n20450 ;
  assign n20452 = n20451 ^ n18955 ;
  assign n20453 = n20452 ^ n18953 ;
  assign n20440 = n20366 ^ n19260 ;
  assign n20441 = ~n20365 & n20440 ;
  assign n20437 = n19494 ^ n19277 ;
  assign n20438 = n20437 ^ n19493 ;
  assign n20439 = n20438 ^ n20366 ;
  assign n20442 = n20441 ^ n20439 ;
  assign n20443 = n20442 ^ n19277 ;
  assign n20444 = n19271 & n20443 ;
  assign n20433 = n20370 ^ n20359 ;
  assign n20434 = n20370 ^ n17988 ;
  assign n20435 = ~n20433 & ~n20434 ;
  assign n20431 = n19277 ^ n18004 ;
  assign n20430 = n17988 ^ x248 ;
  assign n20432 = n20431 ^ n20430 ;
  assign n20436 = n20435 ^ n20432 ;
  assign n20445 = n20444 ^ n20436 ;
  assign n20425 = n20378 ^ n20371 ;
  assign n20428 = ~n20376 & n20425 ;
  assign n20424 = n20376 ^ n20371 ;
  assign n20426 = n20425 ^ n20424 ;
  assign n20427 = x249 & n20426 ;
  assign n20429 = n20428 ^ n20427 ;
  assign n20446 = n20445 ^ n20429 ;
  assign n20421 = n20383 ^ n20379 ;
  assign n20422 = n20380 & ~n20421 ;
  assign n20423 = n20422 ^ n20383 ;
  assign n20447 = n20446 ^ n20423 ;
  assign n20448 = n19114 & ~n20447 ;
  assign n20449 = n20448 ^ n19596 ;
  assign n20454 = n20453 ^ n20449 ;
  assign n20456 = n20454 ^ x395 ;
  assign n20455 = n20454 ^ n20389 ;
  assign n20457 = n20456 ^ n20455 ;
  assign n20458 = n20394 & ~n20457 ;
  assign n20459 = n20458 ^ n20456 ;
  assign n20460 = n20459 ^ x394 ;
  assign n20462 = n20461 ^ n20460 ;
  assign n20465 = n20464 ^ n20462 ;
  assign n20466 = n20465 ^ n19927 ;
  assign n20420 = n18741 & ~n20419 ;
  assign n20467 = n20466 ^ n20420 ;
  assign n20468 = n20467 ^ n18769 ;
  assign n20470 = n20469 ^ n20468 ;
  assign n20496 = n20420 ^ n18769 ;
  assign n20497 = n20467 & n20496 ;
  assign n20498 = n20497 ^ n18769 ;
  assign n20499 = n20498 ^ n19534 ;
  assign n20492 = n20460 & n20461 ;
  assign n20479 = n20446 ^ n19596 ;
  assign n20480 = n20447 & ~n20479 ;
  assign n20481 = n20480 ^ n19596 ;
  assign n20482 = n20481 ^ n19882 ;
  assign n20483 = n19122 & ~n20482 ;
  assign n20484 = n20483 ^ n19591 ;
  assign n20475 = n20452 ^ n20449 ;
  assign n20476 = ~n20453 & n20475 ;
  assign n20477 = n20476 ^ n18953 ;
  assign n20478 = n20477 ^ n18770 ;
  assign n20485 = n20484 ^ n20478 ;
  assign n20487 = n20485 ^ x394 ;
  assign n20486 = n20485 ^ n20454 ;
  assign n20488 = n20487 ^ n20486 ;
  assign n20489 = ~n20459 & n20488 ;
  assign n20490 = n20489 ^ n20487 ;
  assign n20491 = n20490 ^ x393 ;
  assign n20493 = n20492 ^ n20491 ;
  assign n20471 = n19937 ^ n19921 ;
  assign n20472 = n20471 ^ n20464 ;
  assign n20473 = ~n20465 & ~n20472 ;
  assign n20474 = n20473 ^ n20471 ;
  assign n20494 = n20493 ^ n20474 ;
  assign n20495 = n20494 ^ n19967 ;
  assign n20500 = n20499 ^ n20495 ;
  assign n20501 = n20500 ^ x166 ;
  assign n20502 = n20501 ^ n20468 ;
  assign n20503 = n20502 ^ n20500 ;
  assign n20504 = n20470 & ~n20503 ;
  assign n20505 = n20504 ^ n20501 ;
  assign n20530 = n20485 ^ x393 ;
  assign n20531 = ~n20490 & n20530 ;
  assign n20532 = n20531 ^ x393 ;
  assign n20524 = n20484 ^ n20477 ;
  assign n20525 = n20484 ^ n18770 ;
  assign n20526 = n20524 & ~n20525 ;
  assign n20527 = n20526 ^ n18770 ;
  assign n20528 = n20527 ^ n18970 ;
  assign n20519 = n19884 ^ n19882 ;
  assign n20517 = n19697 ^ n19591 ;
  assign n20515 = n19882 ^ n19591 ;
  assign n20516 = n20482 & n20515 ;
  assign n20518 = n20517 ^ n20516 ;
  assign n20520 = n20519 ^ n20518 ;
  assign n20521 = n20520 ^ n19697 ;
  assign n20522 = ~n19130 & n20521 ;
  assign n20523 = n20522 ^ n19697 ;
  assign n20529 = n20528 ^ n20523 ;
  assign n20533 = n20532 ^ n20529 ;
  assign n20534 = n20533 ^ x392 ;
  assign n20514 = ~n20491 & ~n20492 ;
  assign n20535 = n20534 ^ n20514 ;
  assign n20536 = n20535 ^ n20493 ;
  assign n20510 = n19980 ^ n19963 ;
  assign n20511 = n20510 ^ n20493 ;
  assign n20512 = n20510 ^ n20474 ;
  assign n20513 = ~n20511 & n20512 ;
  assign n20537 = n20536 ^ n20513 ;
  assign n20538 = n20537 ^ n20010 ;
  assign n20506 = n20498 ^ n20495 ;
  assign n20507 = ~n20499 & n20506 ;
  assign n20508 = n20507 ^ n19534 ;
  assign n20509 = n20508 ^ n19531 ;
  assign n20539 = n20538 ^ n20509 ;
  assign n20541 = n20539 ^ x165 ;
  assign n20540 = n20539 ^ n20500 ;
  assign n20542 = n20541 ^ n20540 ;
  assign n20543 = ~n20505 & n20542 ;
  assign n20544 = n20543 ^ n20541 ;
  assign n20585 = n20539 ^ x164 ;
  assign n20586 = ~n20544 & n20585 ;
  assign n20587 = n20586 ^ x164 ;
  assign n20565 = n20527 ^ n20523 ;
  assign n20566 = n19886 ^ n19885 ;
  assign n20568 = n20566 ^ n19697 ;
  assign n20567 = n20566 ^ n20519 ;
  assign n20569 = n20568 ^ n20567 ;
  assign n20570 = ~n20518 & ~n20569 ;
  assign n20571 = n20570 ^ n20568 ;
  assign n20572 = ~n19804 & n20571 ;
  assign n20573 = n20572 ^ n19811 ;
  assign n20574 = n20573 ^ n18970 ;
  assign n20575 = n20574 ^ n20573 ;
  assign n20576 = n20575 ^ n20527 ;
  assign n20577 = ~n20565 & n20576 ;
  assign n20578 = n20577 ^ n20574 ;
  assign n20579 = n20578 ^ n18979 ;
  assign n20561 = n20532 ^ x392 ;
  assign n20562 = n20533 & n20561 ;
  assign n20563 = n20562 ^ x392 ;
  assign n20564 = n20563 ^ x407 ;
  assign n20580 = n20579 ^ n20564 ;
  assign n20560 = ~n20514 & ~n20534 ;
  assign n20581 = n20580 ^ n20560 ;
  assign n20555 = n20010 ^ n19982 ;
  assign n20556 = n20555 ^ n20006 ;
  assign n20557 = n20556 ^ n20535 ;
  assign n20558 = n20537 & ~n20557 ;
  assign n20559 = n20558 ^ n20556 ;
  assign n20582 = n20581 ^ n20559 ;
  assign n20583 = n20582 ^ n20051 ;
  assign n20551 = n20538 ^ n20508 ;
  assign n20552 = ~n20509 & ~n20551 ;
  assign n20553 = n20552 ^ n19531 ;
  assign n20554 = n20553 ^ n19527 ;
  assign n20584 = n20583 ^ n20554 ;
  assign n20588 = n20587 ^ n20584 ;
  assign n20602 = n20579 ^ n20563 ;
  assign n20608 = n20566 ^ n19811 ;
  assign n20609 = ~n20571 & ~n20608 ;
  assign n20610 = n20609 ^ n19811 ;
  assign n20607 = n19888 ^ n19887 ;
  assign n20611 = n20610 ^ n20607 ;
  assign n20612 = ~n19840 & ~n20611 ;
  assign n20613 = n20612 ^ n19827 ;
  assign n20603 = n20573 ^ n18979 ;
  assign n20604 = n20578 & n20603 ;
  assign n20605 = n20604 ^ n18979 ;
  assign n20606 = n20605 ^ n18985 ;
  assign n20614 = n20613 ^ n20606 ;
  assign n20615 = n20614 ^ x407 ;
  assign n20616 = n20615 ^ n20579 ;
  assign n20617 = n20616 ^ n20614 ;
  assign n20618 = n20602 & ~n20617 ;
  assign n20619 = n20618 ^ n20615 ;
  assign n20620 = n20619 ^ x406 ;
  assign n20601 = n20560 & ~n20580 ;
  assign n20621 = n20620 ^ n20601 ;
  assign n20595 = n20051 ^ n20024 ;
  assign n20596 = n20595 ^ n20047 ;
  assign n20597 = n20596 ^ n20581 ;
  assign n20598 = n20596 ^ n20559 ;
  assign n20599 = n20597 & ~n20598 ;
  assign n20600 = n20599 ^ n20581 ;
  assign n20622 = n20621 ^ n20600 ;
  assign n20623 = n20622 ^ n20094 ;
  assign n20591 = n20583 ^ n20553 ;
  assign n20592 = n20554 & ~n20591 ;
  assign n20593 = n20592 ^ n19527 ;
  assign n20594 = n20593 ^ n19524 ;
  assign n20624 = n20623 ^ n20594 ;
  assign n20625 = n20624 ^ x163 ;
  assign n20626 = n20625 ^ n20587 ;
  assign n20627 = n20626 ^ n20624 ;
  assign n20628 = ~n20588 & n20627 ;
  assign n20629 = n20628 ^ n20625 ;
  assign n20652 = n19890 ^ n19889 ;
  assign n20650 = n20610 ^ n19846 ;
  assign n20646 = n19840 ^ n19827 ;
  assign n20647 = n20646 ^ n20610 ;
  assign n20648 = n20646 ^ n20607 ;
  assign n20649 = ~n20647 & n20648 ;
  assign n20651 = n20650 ^ n20649 ;
  assign n20653 = n20652 ^ n20651 ;
  assign n20654 = n20653 ^ n19846 ;
  assign n20655 = n19148 & n20654 ;
  assign n20656 = n20655 ^ n19846 ;
  assign n20641 = n20613 ^ n20605 ;
  assign n20642 = n20613 ^ n18985 ;
  assign n20643 = ~n20641 & ~n20642 ;
  assign n20644 = n20643 ^ n18985 ;
  assign n20645 = n20644 ^ n18988 ;
  assign n20657 = n20656 ^ n20645 ;
  assign n20659 = n20657 ^ x406 ;
  assign n20658 = n20657 ^ n20614 ;
  assign n20660 = n20659 ^ n20658 ;
  assign n20661 = n20619 & ~n20660 ;
  assign n20662 = n20661 ^ n20659 ;
  assign n20663 = n20662 ^ x405 ;
  assign n20640 = ~n20601 & n20620 ;
  assign n20664 = n20663 ^ n20640 ;
  assign n20636 = n20107 ^ n20090 ;
  assign n20637 = n20636 ^ n20621 ;
  assign n20638 = n20622 & n20637 ;
  assign n20639 = n20638 ^ n20636 ;
  assign n20665 = n20664 ^ n20639 ;
  assign n20666 = n20665 ^ n20138 ;
  assign n20632 = n20623 ^ n20593 ;
  assign n20633 = n20594 & ~n20632 ;
  assign n20634 = n20633 ^ n19524 ;
  assign n20635 = n20634 ^ n19063 ;
  assign n20667 = n20666 ^ n20635 ;
  assign n20669 = n20667 ^ x162 ;
  assign n20668 = n20667 ^ n20624 ;
  assign n20670 = n20669 ^ n20668 ;
  assign n20671 = ~n20629 & n20670 ;
  assign n20672 = n20671 ^ n20669 ;
  assign n20696 = n19892 ^ n19891 ;
  assign n20692 = n19870 ^ n19846 ;
  assign n20691 = n20652 ^ n19870 ;
  assign n20693 = n20692 ^ n20691 ;
  assign n20694 = n20651 & n20693 ;
  assign n20695 = n20694 ^ n20692 ;
  assign n20697 = n20696 ^ n20695 ;
  assign n20698 = n20697 ^ n19870 ;
  assign n20699 = n19156 & n20698 ;
  assign n20700 = n20699 ^ n19870 ;
  assign n20686 = n20656 ^ n20644 ;
  assign n20687 = n20656 ^ n18988 ;
  assign n20688 = n20686 & ~n20687 ;
  assign n20689 = n20688 ^ n18988 ;
  assign n20690 = n20689 ^ n18991 ;
  assign n20701 = n20700 ^ n20690 ;
  assign n20703 = n20701 ^ x405 ;
  assign n20702 = n20701 ^ n20657 ;
  assign n20704 = n20703 ^ n20702 ;
  assign n20705 = ~n20662 & n20704 ;
  assign n20706 = n20705 ^ n20703 ;
  assign n20707 = n20706 ^ x404 ;
  assign n20685 = ~n20640 & n20663 ;
  assign n20708 = n20707 ^ n20685 ;
  assign n20679 = n20138 ^ n20109 ;
  assign n20680 = n20679 ^ n20134 ;
  assign n20681 = n20680 ^ n20664 ;
  assign n20682 = n20680 ^ n20639 ;
  assign n20683 = ~n20681 & ~n20682 ;
  assign n20684 = n20683 ^ n20664 ;
  assign n20709 = n20708 ^ n20684 ;
  assign n20710 = n20709 ^ n20177 ;
  assign n20675 = n20666 ^ n20634 ;
  assign n20676 = n20635 & n20675 ;
  assign n20677 = n20676 ^ n19063 ;
  assign n20678 = n20677 ^ n19070 ;
  assign n20711 = n20710 ^ n20678 ;
  assign n20713 = n20711 ^ x161 ;
  assign n20712 = n20711 ^ n20667 ;
  assign n20714 = n20713 ^ n20712 ;
  assign n20715 = n20672 & ~n20714 ;
  assign n20716 = n20715 ^ n20713 ;
  assign n20749 = ~n20685 & ~n20707 ;
  assign n20735 = n20696 ^ n19870 ;
  assign n20736 = ~n20695 & ~n20735 ;
  assign n20734 = n19951 ^ n19870 ;
  assign n20737 = n20736 ^ n20734 ;
  assign n20733 = n19894 ^ n19893 ;
  assign n20738 = n20737 ^ n20733 ;
  assign n20739 = n20738 ^ n19951 ;
  assign n20740 = n19164 & n20739 ;
  assign n20741 = n20740 ^ n19951 ;
  assign n20728 = n20700 ^ n20689 ;
  assign n20729 = n20700 ^ n18991 ;
  assign n20730 = ~n20728 & ~n20729 ;
  assign n20731 = n20730 ^ n18991 ;
  assign n20732 = n20731 ^ n18942 ;
  assign n20742 = n20741 ^ n20732 ;
  assign n20744 = n20742 ^ x404 ;
  assign n20743 = n20742 ^ n20701 ;
  assign n20745 = n20744 ^ n20743 ;
  assign n20746 = ~n20706 & n20745 ;
  assign n20747 = n20746 ^ n20744 ;
  assign n20748 = n20747 ^ x403 ;
  assign n20750 = n20749 ^ n20748 ;
  assign n20723 = n20190 ^ n20173 ;
  assign n20724 = n20723 ^ n20708 ;
  assign n20725 = n20723 ^ n20684 ;
  assign n20726 = n20724 & ~n20725 ;
  assign n20727 = n20726 ^ n20708 ;
  assign n20751 = n20750 ^ n20727 ;
  assign n20752 = n20751 ^ n20220 ;
  assign n20719 = n20710 ^ n20677 ;
  assign n20720 = n20678 & ~n20719 ;
  assign n20721 = n20720 ^ n19070 ;
  assign n20722 = n20721 ^ n19079 ;
  assign n20753 = n20752 ^ n20722 ;
  assign n20755 = n20753 ^ x160 ;
  assign n20754 = n20753 ^ n20711 ;
  assign n20756 = n20755 ^ n20754 ;
  assign n20757 = ~n20716 & n20756 ;
  assign n20758 = n20757 ^ n20755 ;
  assign n20791 = n20748 & ~n20749 ;
  assign n20777 = n20733 ^ n19951 ;
  assign n20778 = ~n20737 & ~n20777 ;
  assign n20776 = n19994 ^ n19951 ;
  assign n20779 = n20778 ^ n20776 ;
  assign n20775 = n19896 ^ n19895 ;
  assign n20780 = n20779 ^ n20775 ;
  assign n20781 = n20780 ^ n19994 ;
  assign n20782 = n19172 & n20781 ;
  assign n20783 = n20782 ^ n19994 ;
  assign n20770 = n20741 ^ n20731 ;
  assign n20771 = n20741 ^ n18942 ;
  assign n20772 = ~n20770 & n20771 ;
  assign n20773 = n20772 ^ n18942 ;
  assign n20774 = n20773 ^ n18300 ;
  assign n20784 = n20783 ^ n20774 ;
  assign n20786 = n20784 ^ x403 ;
  assign n20785 = n20784 ^ n20742 ;
  assign n20787 = n20786 ^ n20785 ;
  assign n20788 = ~n20747 & n20787 ;
  assign n20789 = n20788 ^ n20786 ;
  assign n20790 = n20789 ^ x402 ;
  assign n20792 = n20791 ^ n20790 ;
  assign n20765 = n20220 ^ n20192 ;
  assign n20766 = n20765 ^ n20216 ;
  assign n20767 = n20766 ^ n20750 ;
  assign n20768 = ~n20751 & ~n20767 ;
  assign n20769 = n20768 ^ n20766 ;
  assign n20793 = n20792 ^ n20769 ;
  assign n20794 = n20793 ^ n19611 ;
  assign n20761 = n20752 ^ n20721 ;
  assign n20762 = ~n20722 & n20761 ;
  assign n20763 = n20762 ^ n19079 ;
  assign n20764 = n20763 ^ n19087 ;
  assign n20795 = n20794 ^ n20764 ;
  assign n20797 = n20795 ^ x175 ;
  assign n20796 = n20795 ^ n20753 ;
  assign n20798 = n20797 ^ n20796 ;
  assign n20799 = ~n20758 & n20798 ;
  assign n20800 = n20799 ^ n20797 ;
  assign n20833 = n20790 & ~n20791 ;
  assign n20819 = n20775 ^ n19994 ;
  assign n20820 = ~n20779 & ~n20819 ;
  assign n20818 = n20036 ^ n19994 ;
  assign n20821 = n20820 ^ n20818 ;
  assign n20817 = n19898 ^ n19897 ;
  assign n20822 = n20821 ^ n20817 ;
  assign n20823 = n20822 ^ n20036 ;
  assign n20824 = ~n19180 & n20823 ;
  assign n20825 = n20824 ^ n20036 ;
  assign n20812 = n20783 ^ n20773 ;
  assign n20813 = n20783 ^ n18300 ;
  assign n20814 = n20812 & ~n20813 ;
  assign n20815 = n20814 ^ n18300 ;
  assign n20816 = n20815 ^ n18448 ;
  assign n20826 = n20825 ^ n20816 ;
  assign n20828 = n20826 ^ x402 ;
  assign n20827 = n20826 ^ n20784 ;
  assign n20829 = n20828 ^ n20827 ;
  assign n20830 = n20789 & ~n20829 ;
  assign n20831 = n20830 ^ n20828 ;
  assign n20832 = n20831 ^ x401 ;
  assign n20834 = n20833 ^ n20832 ;
  assign n20807 = n20234 ^ n19611 ;
  assign n20808 = n20807 ^ n20258 ;
  assign n20809 = n20808 ^ n20792 ;
  assign n20810 = ~n20793 & n20809 ;
  assign n20811 = n20810 ^ n20808 ;
  assign n20835 = n20834 ^ n20811 ;
  assign n20836 = n20835 ^ n19606 ;
  assign n20803 = n20794 ^ n20763 ;
  assign n20804 = n20764 & ~n20803 ;
  assign n20805 = n20804 ^ n19087 ;
  assign n20806 = n20805 ^ n18928 ;
  assign n20837 = n20836 ^ n20806 ;
  assign n20839 = n20837 ^ x174 ;
  assign n20838 = n20837 ^ n20795 ;
  assign n20840 = n20839 ^ n20838 ;
  assign n20841 = n20800 & ~n20840 ;
  assign n20842 = n20841 ^ n20839 ;
  assign n20876 = ~n20832 & ~n20833 ;
  assign n20864 = n20825 ^ n20815 ;
  assign n20865 = n20825 ^ n18448 ;
  assign n20866 = ~n20864 & ~n20865 ;
  assign n20867 = n20866 ^ n18448 ;
  assign n20868 = n20867 ^ n18462 ;
  assign n20859 = n19900 ^ n19899 ;
  assign n20854 = n20073 ^ n20036 ;
  assign n20855 = n20854 ^ n20073 ;
  assign n20856 = n20855 ^ n20817 ;
  assign n20857 = ~n20821 & ~n20856 ;
  assign n20858 = n20857 ^ n20854 ;
  assign n20860 = n20859 ^ n20858 ;
  assign n20861 = n20860 ^ n20073 ;
  assign n20862 = n19187 & ~n20861 ;
  assign n20863 = n20862 ^ n20073 ;
  assign n20869 = n20868 ^ n20863 ;
  assign n20871 = n20869 ^ x401 ;
  assign n20870 = n20869 ^ n20826 ;
  assign n20872 = n20871 ^ n20870 ;
  assign n20873 = n20831 & ~n20872 ;
  assign n20874 = n20873 ^ n20871 ;
  assign n20875 = n20874 ^ x400 ;
  assign n20877 = n20876 ^ n20875 ;
  assign n20849 = n20314 ^ n20297 ;
  assign n20850 = n20849 ^ n20834 ;
  assign n20851 = n20849 ^ n20811 ;
  assign n20852 = ~n20850 & n20851 ;
  assign n20853 = n20852 ^ n20834 ;
  assign n20878 = n20877 ^ n20853 ;
  assign n20879 = n20878 ^ n19601 ;
  assign n20845 = n20836 ^ n20805 ;
  assign n20846 = ~n20806 & n20845 ;
  assign n20847 = n20846 ^ n18928 ;
  assign n20848 = n20847 ^ n18902 ;
  assign n20880 = n20879 ^ n20848 ;
  assign n20882 = n20880 ^ x173 ;
  assign n20881 = n20880 ^ n20837 ;
  assign n20883 = n20882 ^ n20881 ;
  assign n20884 = n20842 & ~n20883 ;
  assign n20885 = n20884 ^ n20882 ;
  assign n20916 = n20875 & n20876 ;
  assign n20911 = n20869 ^ x400 ;
  assign n20912 = ~n20874 & n20911 ;
  assign n20913 = n20912 ^ x400 ;
  assign n20914 = n20913 ^ x415 ;
  assign n20896 = n20867 ^ n20863 ;
  assign n20897 = n19902 ^ n19901 ;
  assign n20899 = n20897 ^ n20073 ;
  assign n20898 = n20897 ^ n20859 ;
  assign n20900 = n20899 ^ n20898 ;
  assign n20901 = ~n20858 & n20900 ;
  assign n20902 = n20901 ^ n20899 ;
  assign n20903 = ~n20115 & ~n20902 ;
  assign n20904 = n20903 ^ n20122 ;
  assign n20905 = n20904 ^ n18462 ;
  assign n20906 = n20905 ^ n20904 ;
  assign n20907 = n20906 ^ n20867 ;
  assign n20908 = ~n20896 & ~n20907 ;
  assign n20909 = n20908 ^ n20905 ;
  assign n20910 = n20909 ^ n19022 ;
  assign n20915 = n20914 ^ n20910 ;
  assign n20917 = n20916 ^ n20915 ;
  assign n20892 = n20353 ^ n20316 ;
  assign n20893 = n20892 ^ n20877 ;
  assign n20894 = ~n20878 & n20893 ;
  assign n20895 = n20894 ^ n20892 ;
  assign n20918 = n20917 ^ n20895 ;
  assign n20919 = n20918 ^ n20383 ;
  assign n20888 = n20879 ^ n20847 ;
  assign n20889 = ~n20848 & n20888 ;
  assign n20890 = n20889 ^ n18902 ;
  assign n20891 = n20890 ^ n19577 ;
  assign n20920 = n20919 ^ n20891 ;
  assign n20922 = n20920 ^ x172 ;
  assign n20921 = n20920 ^ n20880 ;
  assign n20923 = n20922 ^ n20921 ;
  assign n20924 = ~n20885 & n20923 ;
  assign n20925 = n20924 ^ n20922 ;
  assign n20926 = n20925 ^ x171 ;
  assign n20545 = n20544 ^ x164 ;
  assign n20546 = n20469 ^ x166 ;
  assign n20547 = n20546 ^ n20468 ;
  assign n20548 = n20505 ^ x165 ;
  assign n20549 = ~n20547 & n20548 ;
  assign n20550 = n20545 & n20549 ;
  assign n20589 = n20588 ^ x163 ;
  assign n20590 = n20550 & n20589 ;
  assign n20630 = n20629 ^ x162 ;
  assign n20631 = n20590 & n20630 ;
  assign n20673 = n20672 ^ x161 ;
  assign n20674 = ~n20631 & n20673 ;
  assign n20717 = n20716 ^ x160 ;
  assign n20718 = ~n20674 & n20717 ;
  assign n20759 = n20758 ^ x175 ;
  assign n20760 = ~n20718 & ~n20759 ;
  assign n20801 = n20800 ^ x174 ;
  assign n20802 = ~n20760 & ~n20801 ;
  assign n20843 = n20842 ^ x173 ;
  assign n20844 = n20802 & ~n20843 ;
  assign n20886 = n20885 ^ x172 ;
  assign n20887 = ~n20844 & ~n20886 ;
  assign n21814 = n20926 ^ n20887 ;
  assign n21651 = n20808 ^ n20769 ;
  assign n21652 = n21651 ^ n20792 ;
  assign n21626 = n20766 ^ n20727 ;
  assign n21627 = n21626 ^ n20750 ;
  assign n21653 = n21652 ^ n21627 ;
  assign n21631 = n20589 ^ n20550 ;
  assign n21414 = n20472 ^ n20462 ;
  assign n21293 = n20400 ^ n20399 ;
  assign n21231 = n19934 ^ x391 ;
  assign n21232 = n21231 ^ n20697 ;
  assign n21099 = n20571 ^ n19811 ;
  assign n20942 = n20913 ^ n20910 ;
  assign n20948 = n20897 ^ n20122 ;
  assign n20949 = n20902 & ~n20948 ;
  assign n20950 = n20949 ^ n20122 ;
  assign n20947 = n19904 ^ n19903 ;
  assign n20951 = n20950 ^ n20947 ;
  assign n20952 = ~n19199 & n20951 ;
  assign n20953 = n20952 ^ n20162 ;
  assign n20943 = n20904 ^ n19022 ;
  assign n20944 = n20909 & ~n20943 ;
  assign n20945 = n20944 ^ n19022 ;
  assign n20946 = n20945 ^ n18934 ;
  assign n20954 = n20953 ^ n20946 ;
  assign n20955 = n20954 ^ x415 ;
  assign n20956 = n20955 ^ n20910 ;
  assign n20957 = n20956 ^ n20954 ;
  assign n20958 = n20942 & ~n20957 ;
  assign n20959 = n20958 ^ n20955 ;
  assign n20988 = n19906 ^ n19905 ;
  assign n20986 = n20947 ^ n20204 ;
  assign n20983 = n20162 ^ n19199 ;
  assign n20984 = n20983 ^ n20947 ;
  assign n20985 = ~n20951 & ~n20984 ;
  assign n20987 = n20986 ^ n20985 ;
  assign n20989 = n20988 ^ n20987 ;
  assign n20990 = n20989 ^ n20204 ;
  assign n20991 = ~n19030 & n20990 ;
  assign n20992 = n20991 ^ n20204 ;
  assign n20978 = n20953 ^ n20945 ;
  assign n20979 = n20953 ^ n18934 ;
  assign n20980 = ~n20978 & n20979 ;
  assign n20981 = n20980 ^ n18934 ;
  assign n20982 = n20981 ^ n18652 ;
  assign n20993 = n20992 ^ n20982 ;
  assign n20995 = n20993 ^ x414 ;
  assign n20994 = n20993 ^ n20954 ;
  assign n20996 = n20995 ^ n20994 ;
  assign n20997 = ~n20959 & n20996 ;
  assign n20998 = n20997 ^ n20995 ;
  assign n21030 = n19909 ^ n19907 ;
  assign n21026 = n20246 ^ n20204 ;
  assign n21025 = n20988 ^ n20246 ;
  assign n21027 = n21026 ^ n21025 ;
  assign n21028 = n20987 & n21027 ;
  assign n21029 = n21028 ^ n21026 ;
  assign n21031 = n21030 ^ n21029 ;
  assign n21032 = n21031 ^ n20246 ;
  assign n21033 = n19221 & n21032 ;
  assign n21034 = n21033 ^ n20246 ;
  assign n21020 = n20992 ^ n20981 ;
  assign n21021 = n20992 ^ n18652 ;
  assign n21022 = ~n21020 & ~n21021 ;
  assign n21023 = n21022 ^ n18652 ;
  assign n21024 = n21023 ^ n18673 ;
  assign n21035 = n21034 ^ n21024 ;
  assign n21037 = n21035 ^ x413 ;
  assign n21036 = n21035 ^ n20993 ;
  assign n21038 = n21037 ^ n21036 ;
  assign n21039 = n20998 & ~n21038 ;
  assign n21040 = n21039 ^ n21037 ;
  assign n21041 = n21040 ^ x412 ;
  assign n20999 = n20998 ^ x413 ;
  assign n20960 = n20959 ^ x414 ;
  assign n20961 = n20915 & ~n20916 ;
  assign n21000 = n20960 & ~n20961 ;
  assign n21042 = n20999 & ~n21000 ;
  assign n21082 = ~n21041 & n21042 ;
  assign n21070 = n19911 ^ n19910 ;
  assign n21066 = n20285 ^ n20246 ;
  assign n21065 = n21030 ^ n20285 ;
  assign n21067 = n21066 ^ n21065 ;
  assign n21068 = ~n21029 & ~n21067 ;
  assign n21069 = n21068 ^ n21066 ;
  assign n21071 = n21070 ^ n21069 ;
  assign n21072 = n21071 ^ n20285 ;
  assign n21073 = n20278 & n21072 ;
  assign n21074 = n21073 ^ n20285 ;
  assign n21060 = n21034 ^ n21023 ;
  assign n21061 = n21034 ^ n18673 ;
  assign n21062 = ~n21060 & ~n21061 ;
  assign n21063 = n21062 ^ n18673 ;
  assign n21064 = n21063 ^ n18756 ;
  assign n21075 = n21074 ^ n21064 ;
  assign n21077 = n21075 ^ x412 ;
  assign n21076 = n21075 ^ n21035 ;
  assign n21078 = n21077 ^ n21076 ;
  assign n21079 = ~n21040 & n21078 ;
  assign n21080 = n21079 ^ n21077 ;
  assign n21081 = n21080 ^ x411 ;
  assign n21083 = n21082 ^ n21081 ;
  assign n21100 = n21099 ^ n21083 ;
  assign n21123 = ~n21081 & ~n21082 ;
  assign n21111 = n19913 ^ n19912 ;
  assign n21107 = n20327 ^ n20285 ;
  assign n21106 = n21070 ^ n20327 ;
  assign n21108 = n21107 ^ n21106 ;
  assign n21109 = ~n21069 & ~n21108 ;
  assign n21110 = n21109 ^ n21107 ;
  assign n21112 = n21111 ^ n21110 ;
  assign n21113 = n21112 ^ n20327 ;
  assign n21114 = ~n19247 & n21113 ;
  assign n21115 = n21114 ^ n20327 ;
  assign n21101 = n21074 ^ n21063 ;
  assign n21102 = n21074 ^ n18756 ;
  assign n21103 = ~n21101 & ~n21102 ;
  assign n21104 = n21103 ^ n18756 ;
  assign n21105 = n21104 ^ n19240 ;
  assign n21116 = n21115 ^ n21105 ;
  assign n21118 = n21116 ^ x411 ;
  assign n21117 = n21116 ^ n21075 ;
  assign n21119 = n21118 ^ n21117 ;
  assign n21120 = n21080 & ~n21119 ;
  assign n21121 = n21120 ^ n21118 ;
  assign n21122 = n21121 ^ x410 ;
  assign n21124 = n21123 ^ n21122 ;
  assign n21043 = n21042 ^ n21041 ;
  assign n21001 = n21000 ^ n20999 ;
  assign n21044 = n21043 ^ n21001 ;
  assign n21016 = n20515 ^ n20481 ;
  assign n21017 = n21016 ^ n21001 ;
  assign n20962 = n20961 ^ n20960 ;
  assign n20936 = n20383 ^ n20355 ;
  assign n20937 = n20936 ^ n20379 ;
  assign n20938 = n20937 ^ n20917 ;
  assign n20939 = n20937 ^ n20895 ;
  assign n20940 = n20938 & ~n20939 ;
  assign n20941 = n20940 ^ n20917 ;
  assign n20963 = n20962 ^ n20941 ;
  assign n20973 = n20423 ^ n19596 ;
  assign n20974 = n20973 ^ n20446 ;
  assign n20975 = n20974 ^ n20962 ;
  assign n20976 = n20963 & ~n20975 ;
  assign n20977 = n20976 ^ n20974 ;
  assign n21018 = n21016 ^ n20977 ;
  assign n21019 = ~n21017 & n21018 ;
  assign n21045 = n21044 ^ n21019 ;
  assign n21084 = n21043 ^ n20520 ;
  assign n21085 = ~n21045 & ~n21084 ;
  assign n21086 = n21085 ^ n20520 ;
  assign n21125 = n21124 ^ n21086 ;
  assign n21126 = n21125 ^ n21083 ;
  assign n21127 = n21126 ^ n21124 ;
  assign n21128 = ~n21100 & ~n21127 ;
  assign n21129 = n21128 ^ n21125 ;
  assign n21171 = n20646 ^ n20611 ;
  assign n21172 = n21171 ^ n21124 ;
  assign n21173 = n21129 & n21172 ;
  assign n21168 = ~n21122 & n21123 ;
  assign n21156 = n19916 ^ n19914 ;
  assign n21152 = n20367 ^ n20327 ;
  assign n21151 = n21111 ^ n20367 ;
  assign n21153 = n21152 ^ n21151 ;
  assign n21154 = ~n21110 & ~n21153 ;
  assign n21155 = n21154 ^ n21152 ;
  assign n21157 = n21156 ^ n21155 ;
  assign n21158 = n21157 ^ n20367 ;
  assign n21159 = ~n19260 & ~n21158 ;
  assign n21160 = n21159 ^ n20367 ;
  assign n21146 = n21115 ^ n21104 ;
  assign n21147 = n21115 ^ n19240 ;
  assign n21148 = ~n21146 & n21147 ;
  assign n21149 = n21148 ^ n19240 ;
  assign n21150 = n21149 ^ n18813 ;
  assign n21161 = n21160 ^ n21150 ;
  assign n21163 = n21161 ^ x410 ;
  assign n21162 = n21161 ^ n21116 ;
  assign n21164 = n21163 ^ n21162 ;
  assign n21165 = n21121 & ~n21164 ;
  assign n21166 = n21165 ^ n21163 ;
  assign n21167 = n21166 ^ x409 ;
  assign n21169 = n21168 ^ n21167 ;
  assign n21170 = n21169 ^ n21124 ;
  assign n21174 = n21173 ^ n21170 ;
  assign n21208 = n21169 ^ n20653 ;
  assign n21209 = n21174 & n21208 ;
  assign n21210 = n21209 ^ n20653 ;
  assign n21204 = n21168 ^ n21161 ;
  assign n21205 = ~n21166 & ~n21204 ;
  assign n21202 = n21168 ^ n21166 ;
  assign n21203 = ~x409 & n21202 ;
  assign n21206 = n21205 ^ n21203 ;
  assign n21196 = n21156 ^ n20367 ;
  assign n21197 = ~n21155 & ~n21196 ;
  assign n21193 = n20442 ^ n19917 ;
  assign n21194 = n21193 ^ n19918 ;
  assign n21195 = n21194 ^ n21156 ;
  assign n21198 = n21197 ^ n21195 ;
  assign n21199 = n21198 ^ n20442 ;
  assign n21200 = ~n19277 & n21199 ;
  assign n21190 = n20442 ^ n19271 ;
  assign n21189 = n18813 ^ x408 ;
  assign n21191 = n21190 ^ n21189 ;
  assign n21186 = n21160 ^ n21149 ;
  assign n21187 = n21160 ^ n18813 ;
  assign n21188 = ~n21186 & ~n21187 ;
  assign n21192 = n21191 ^ n21188 ;
  assign n21201 = n21200 ^ n21192 ;
  assign n21207 = n21206 ^ n21201 ;
  assign n21211 = n21210 ^ n21207 ;
  assign n21229 = n21210 ^ n20697 ;
  assign n21230 = n21211 & ~n21229 ;
  assign n21233 = n21232 ^ n21230 ;
  assign n21248 = n21231 ^ n20738 ;
  assign n21249 = ~n21233 & n21248 ;
  assign n21250 = n21249 ^ n21231 ;
  assign n21266 = n21250 ^ n20780 ;
  assign n21267 = n20822 ^ n20397 ;
  assign n21268 = n21267 ^ n20822 ;
  assign n21269 = n21268 ^ n21250 ;
  assign n21270 = n21266 & n21269 ;
  assign n21271 = n21270 ^ n21267 ;
  assign n21289 = n20860 ^ n20822 ;
  assign n21272 = n20398 ^ n20397 ;
  assign n21288 = n21272 ^ n20860 ;
  assign n21290 = n21289 ^ n21288 ;
  assign n21291 = n21271 & ~n21290 ;
  assign n21292 = n21291 ^ n21289 ;
  assign n21294 = n21293 ^ n21292 ;
  assign n21295 = n21294 ^ n20860 ;
  assign n21296 = n21295 ^ n20073 ;
  assign n21273 = n21272 ^ n21271 ;
  assign n21274 = n21273 ^ n20822 ;
  assign n21275 = n21274 ^ n20036 ;
  assign n21283 = n21275 ^ n19180 ;
  assign n21251 = n21250 ^ n20397 ;
  assign n21252 = n21251 ^ n19994 ;
  assign n21234 = n21233 ^ n19951 ;
  assign n21243 = n21234 ^ n19164 ;
  assign n21175 = n21174 ^ n19846 ;
  assign n21176 = n21175 ^ n19840 ;
  assign n21046 = n21045 ^ n19697 ;
  assign n20932 = n20919 ^ n20890 ;
  assign n20933 = n20891 & ~n20932 ;
  assign n20934 = n20933 ^ n19577 ;
  assign n20935 = n20934 ^ n19114 ;
  assign n20964 = n20963 ^ n19596 ;
  assign n20969 = n20964 ^ n20934 ;
  assign n20970 = ~n20935 & n20969 ;
  assign n20971 = n20970 ^ n19114 ;
  assign n20972 = n20971 ^ n19122 ;
  assign n21002 = n21001 ^ n20977 ;
  assign n21003 = n21002 ^ n19591 ;
  assign n21012 = n21003 ^ n20971 ;
  assign n21013 = n20972 & ~n21012 ;
  assign n21014 = n21013 ^ n19122 ;
  assign n21059 = n21046 ^ n21014 ;
  assign n21087 = n21086 ^ n21083 ;
  assign n21088 = n21087 ^ n19811 ;
  assign n21089 = n21088 ^ n19130 ;
  assign n21090 = n21089 ^ n21046 ;
  assign n21091 = n21090 ^ n21088 ;
  assign n21092 = n21059 & n21091 ;
  assign n21093 = n21092 ^ n21089 ;
  assign n21131 = n20646 ^ n19804 ;
  assign n21132 = n21131 ^ n21129 ;
  assign n21098 = n21088 ^ n20646 ;
  assign n21130 = n21129 ^ n21098 ;
  assign n21133 = n21132 ^ n21130 ;
  assign n21134 = ~n21093 & n21133 ;
  assign n21135 = n21134 ^ n21132 ;
  assign n21144 = n21129 ^ n19827 ;
  assign n21145 = ~n21135 & n21144 ;
  assign n21177 = n21176 ^ n21145 ;
  assign n21213 = n21175 ^ n19148 ;
  assign n21214 = ~n21177 & ~n21213 ;
  assign n21215 = n21214 ^ n19148 ;
  assign n21216 = n21215 ^ n19156 ;
  assign n21212 = n21211 ^ n19870 ;
  assign n21225 = n21215 ^ n21212 ;
  assign n21226 = n21216 & ~n21225 ;
  assign n21227 = n21226 ^ n19156 ;
  assign n21244 = n21234 ^ n21227 ;
  assign n21245 = ~n21243 & n21244 ;
  assign n21246 = n21245 ^ n19164 ;
  assign n21261 = n21252 ^ n21246 ;
  assign n21262 = n21252 ^ n19172 ;
  assign n21263 = n21261 & ~n21262 ;
  assign n21264 = n21263 ^ n19172 ;
  assign n21284 = n21275 ^ n21264 ;
  assign n21285 = n21283 & n21284 ;
  assign n21286 = n21285 ^ n19180 ;
  assign n21309 = n21296 ^ n21286 ;
  assign n21313 = n21293 ^ n20860 ;
  assign n21314 = n21292 & n21313 ;
  assign n21315 = n21314 ^ n20860 ;
  assign n21311 = n20402 ^ n20401 ;
  assign n21310 = n20902 ^ n20122 ;
  assign n21312 = n21311 ^ n21310 ;
  assign n21316 = n21315 ^ n21312 ;
  assign n21317 = n21316 ^ n21310 ;
  assign n21318 = n21317 ^ n20122 ;
  assign n21319 = n21318 ^ n19187 ;
  assign n21320 = n21319 ^ n21286 ;
  assign n21321 = n21320 ^ n21318 ;
  assign n21322 = ~n21309 & ~n21321 ;
  assign n21323 = n21322 ^ n21319 ;
  assign n21324 = n21323 ^ n20115 ;
  assign n21094 = n21093 ^ n19804 ;
  assign n20965 = n20964 ^ n20935 ;
  assign n20928 = n20920 ^ x171 ;
  assign n20929 = n20925 & ~n20928 ;
  assign n20930 = n20929 ^ x171 ;
  assign n20968 = n20965 ^ n20930 ;
  assign n21004 = n21003 ^ n20972 ;
  assign n21005 = n21004 ^ x170 ;
  assign n21006 = n21005 ^ n20965 ;
  assign n21007 = n21006 ^ n21004 ;
  assign n21008 = n20968 & ~n21007 ;
  assign n21009 = n21008 ^ n21005 ;
  assign n21015 = n21014 ^ n19130 ;
  assign n21047 = n21046 ^ n21015 ;
  assign n21049 = n21047 ^ x169 ;
  assign n21048 = n21047 ^ n21004 ;
  assign n21050 = n21049 ^ n21048 ;
  assign n21051 = ~n21009 & n21050 ;
  assign n21052 = n21051 ^ n21049 ;
  assign n21055 = n21047 ^ x168 ;
  assign n21056 = ~n21052 & n21055 ;
  assign n21057 = n21056 ^ x168 ;
  assign n21097 = n21094 ^ n21057 ;
  assign n21136 = n21135 ^ n19840 ;
  assign n21137 = n21136 ^ x183 ;
  assign n21138 = n21137 ^ n21094 ;
  assign n21139 = n21138 ^ n21136 ;
  assign n21140 = n21097 & ~n21139 ;
  assign n21141 = n21140 ^ n21137 ;
  assign n21178 = n21177 ^ n19148 ;
  assign n21180 = n21178 ^ x182 ;
  assign n21179 = n21178 ^ n21136 ;
  assign n21181 = n21180 ^ n21179 ;
  assign n21182 = n21141 & ~n21181 ;
  assign n21183 = n21182 ^ n21180 ;
  assign n21217 = n21216 ^ n21212 ;
  assign n21219 = n21217 ^ x181 ;
  assign n21218 = n21217 ^ n21178 ;
  assign n21220 = n21219 ^ n21218 ;
  assign n21221 = ~n21183 & n21220 ;
  assign n21222 = n21221 ^ n21219 ;
  assign n21228 = n21227 ^ n19164 ;
  assign n21235 = n21234 ^ n21228 ;
  assign n21237 = n21235 ^ x180 ;
  assign n21236 = n21235 ^ n21217 ;
  assign n21238 = n21237 ^ n21236 ;
  assign n21239 = ~n21222 & n21238 ;
  assign n21240 = n21239 ^ n21237 ;
  assign n21247 = n21246 ^ n19172 ;
  assign n21253 = n21252 ^ n21247 ;
  assign n21255 = n21253 ^ x179 ;
  assign n21254 = n21253 ^ n21235 ;
  assign n21256 = n21255 ^ n21254 ;
  assign n21257 = n21240 & ~n21256 ;
  assign n21258 = n21257 ^ n21255 ;
  assign n21277 = n21253 ^ x178 ;
  assign n21278 = n21258 & ~n21277 ;
  assign n21279 = n21278 ^ x178 ;
  assign n21265 = n21264 ^ n19180 ;
  assign n21276 = n21275 ^ n21265 ;
  assign n21280 = n21279 ^ n21276 ;
  assign n21287 = n21286 ^ n19187 ;
  assign n21297 = n21296 ^ n21287 ;
  assign n21299 = n21297 ^ x177 ;
  assign n21298 = n21297 ^ n21279 ;
  assign n21300 = n21299 ^ n21298 ;
  assign n21301 = ~n21280 & n21300 ;
  assign n21302 = n21301 ^ n21299 ;
  assign n21305 = n21297 ^ x176 ;
  assign n21306 = ~n21302 & n21305 ;
  assign n21307 = n21306 ^ x176 ;
  assign n21327 = n21324 ^ n21307 ;
  assign n21335 = n20983 ^ n20115 ;
  assign n21332 = n20404 ^ n20403 ;
  assign n21329 = n21315 ^ n21311 ;
  assign n21330 = n21312 & ~n21329 ;
  assign n21331 = n21330 ^ n21315 ;
  assign n21333 = n21332 ^ n21331 ;
  assign n21336 = n21335 ^ n21333 ;
  assign n21328 = n21318 ^ n20983 ;
  assign n21334 = n21333 ^ n21328 ;
  assign n21337 = n21336 ^ n21334 ;
  assign n21338 = ~n21323 & ~n21337 ;
  assign n21339 = n21338 ^ n21336 ;
  assign n21340 = n21339 ^ n19199 ;
  assign n21341 = n21340 ^ x191 ;
  assign n21342 = n21341 ^ n21307 ;
  assign n21343 = n21342 ^ n21340 ;
  assign n21344 = n21327 & n21343 ;
  assign n21345 = n21344 ^ n21341 ;
  assign n21358 = n21333 ^ n20162 ;
  assign n21359 = ~n21339 & n21358 ;
  assign n21348 = n20983 ^ n20951 ;
  assign n21349 = n21348 ^ n21331 ;
  assign n21350 = n20406 ^ n20405 ;
  assign n21351 = n21350 ^ n21332 ;
  assign n21352 = n21351 ^ n21350 ;
  assign n21353 = n21352 ^ n21331 ;
  assign n21354 = ~n21349 & n21353 ;
  assign n21355 = n21354 ^ n21351 ;
  assign n21356 = n21355 ^ n20204 ;
  assign n21357 = n21356 ^ n19199 ;
  assign n21360 = n21359 ^ n21357 ;
  assign n21361 = n21360 ^ n19030 ;
  assign n21363 = n21361 ^ x190 ;
  assign n21362 = n21361 ^ n21340 ;
  assign n21364 = n21363 ^ n21362 ;
  assign n21365 = n21345 & ~n21364 ;
  assign n21366 = n21365 ^ n21363 ;
  assign n21378 = n20408 ^ n20407 ;
  assign n21374 = n21031 ^ n20989 ;
  assign n21373 = n21350 ^ n21031 ;
  assign n21375 = n21374 ^ n21373 ;
  assign n21376 = n21355 & ~n21375 ;
  assign n21377 = n21376 ^ n21374 ;
  assign n21379 = n21378 ^ n21377 ;
  assign n21380 = n21379 ^ n21031 ;
  assign n21381 = n21380 ^ n20246 ;
  assign n21369 = n21356 ^ n19030 ;
  assign n21370 = ~n21360 & n21369 ;
  assign n21371 = n21370 ^ n19030 ;
  assign n21372 = n21371 ^ n19221 ;
  assign n21382 = n21381 ^ n21372 ;
  assign n21384 = n21382 ^ x189 ;
  assign n21383 = n21382 ^ n21361 ;
  assign n21385 = n21384 ^ n21383 ;
  assign n21386 = n21366 & ~n21385 ;
  assign n21387 = n21386 ^ n21384 ;
  assign n21400 = n20410 ^ n20409 ;
  assign n21396 = n21071 ^ n21031 ;
  assign n21395 = n21378 ^ n21071 ;
  assign n21397 = n21396 ^ n21395 ;
  assign n21398 = ~n21377 & ~n21397 ;
  assign n21399 = n21398 ^ n21396 ;
  assign n21401 = n21400 ^ n21399 ;
  assign n21402 = n21401 ^ n21071 ;
  assign n21403 = n21402 ^ n20285 ;
  assign n21390 = n21381 ^ n21371 ;
  assign n21391 = n21381 ^ n19221 ;
  assign n21392 = ~n21390 & ~n21391 ;
  assign n21393 = n21392 ^ n19221 ;
  assign n21394 = n21393 ^ n20278 ;
  assign n21404 = n21403 ^ n21394 ;
  assign n21406 = n21404 ^ x188 ;
  assign n21405 = n21404 ^ n21382 ;
  assign n21407 = n21406 ^ n21405 ;
  assign n21408 = ~n21387 & n21407 ;
  assign n21409 = n21408 ^ n21406 ;
  assign n21410 = n21409 ^ x187 ;
  assign n20927 = n20887 & n20926 ;
  assign n20931 = n20930 ^ x170 ;
  assign n20966 = n20965 ^ n20931 ;
  assign n20967 = n20927 & n20966 ;
  assign n21010 = n21009 ^ x169 ;
  assign n21011 = ~n20967 & n21010 ;
  assign n21053 = n21052 ^ x168 ;
  assign n21054 = n21011 & n21053 ;
  assign n21058 = n21057 ^ x183 ;
  assign n21095 = n21094 ^ n21058 ;
  assign n21096 = n21054 & ~n21095 ;
  assign n21142 = n21141 ^ x182 ;
  assign n21143 = ~n21096 & n21142 ;
  assign n21184 = n21183 ^ x181 ;
  assign n21185 = ~n21143 & n21184 ;
  assign n21223 = n21222 ^ x180 ;
  assign n21224 = ~n21185 & ~n21223 ;
  assign n21241 = n21240 ^ x179 ;
  assign n21242 = n21224 & n21241 ;
  assign n21259 = n21258 ^ x178 ;
  assign n21260 = n21242 & n21259 ;
  assign n21281 = n21280 ^ x177 ;
  assign n21282 = n21260 & ~n21281 ;
  assign n21303 = n21302 ^ x176 ;
  assign n21304 = n21282 & ~n21303 ;
  assign n21308 = n21307 ^ x191 ;
  assign n21325 = n21324 ^ n21308 ;
  assign n21326 = n21304 & n21325 ;
  assign n21346 = n21345 ^ x190 ;
  assign n21347 = n21326 & n21346 ;
  assign n21367 = n21366 ^ x189 ;
  assign n21368 = n21347 & n21367 ;
  assign n21388 = n21387 ^ x188 ;
  assign n21389 = n21368 & ~n21388 ;
  assign n21411 = n21410 ^ n21389 ;
  assign n21412 = n20463 ^ n20418 ;
  assign n21413 = ~n21411 & n21412 ;
  assign n21415 = n21414 ^ n21413 ;
  assign n21428 = n20412 ^ n20411 ;
  assign n21424 = n21112 ^ n21071 ;
  assign n21423 = n21400 ^ n21112 ;
  assign n21425 = n21424 ^ n21423 ;
  assign n21426 = ~n21399 & n21425 ;
  assign n21427 = n21426 ^ n21424 ;
  assign n21429 = n21428 ^ n21427 ;
  assign n21430 = n21429 ^ n21112 ;
  assign n21431 = n21430 ^ n20327 ;
  assign n21418 = n21403 ^ n21393 ;
  assign n21419 = n21403 ^ n20278 ;
  assign n21420 = n21418 & ~n21419 ;
  assign n21421 = n21420 ^ n20278 ;
  assign n21422 = n21421 ^ n19247 ;
  assign n21432 = n21431 ^ n21422 ;
  assign n21434 = n21432 ^ x187 ;
  assign n21433 = n21432 ^ n21404 ;
  assign n21435 = n21434 ^ n21433 ;
  assign n21436 = n21409 & ~n21435 ;
  assign n21437 = n21436 ^ n21434 ;
  assign n21438 = n21437 ^ x186 ;
  assign n21417 = n21389 & n21410 ;
  assign n21439 = n21438 ^ n21417 ;
  assign n21416 = n20512 ^ n20493 ;
  assign n21440 = n21439 ^ n21416 ;
  assign n21441 = n21440 ^ n21413 ;
  assign n21442 = n21441 ^ n21416 ;
  assign n21443 = n21415 & n21442 ;
  assign n21444 = n21443 ^ n21440 ;
  assign n21458 = n20414 ^ n20413 ;
  assign n21454 = n21157 ^ n21112 ;
  assign n21453 = n21428 ^ n21157 ;
  assign n21455 = n21454 ^ n21453 ;
  assign n21456 = ~n21427 & ~n21455 ;
  assign n21457 = n21456 ^ n21454 ;
  assign n21459 = n21458 ^ n21457 ;
  assign n21460 = n21459 ^ n21157 ;
  assign n21461 = n21460 ^ n20367 ;
  assign n21448 = n21431 ^ n21421 ;
  assign n21449 = n21431 ^ n19247 ;
  assign n21450 = n21448 & n21449 ;
  assign n21451 = n21450 ^ n19247 ;
  assign n21452 = n21451 ^ n19260 ;
  assign n21462 = n21461 ^ n21452 ;
  assign n21464 = n21462 ^ x186 ;
  assign n21463 = n21462 ^ n21432 ;
  assign n21465 = n21464 ^ n21463 ;
  assign n21466 = ~n21437 & n21465 ;
  assign n21467 = n21466 ^ n21464 ;
  assign n21468 = n21467 ^ x185 ;
  assign n21447 = n21417 & ~n21438 ;
  assign n21469 = n21468 ^ n21447 ;
  assign n21445 = n20556 ^ n20537 ;
  assign n21470 = n21469 ^ n21445 ;
  assign n21446 = n21445 ^ n21416 ;
  assign n21471 = n21470 ^ n21446 ;
  assign n21472 = n21444 & ~n21471 ;
  assign n21473 = n21472 ^ n21446 ;
  assign n21492 = n21462 ^ n21447 ;
  assign n21495 = n21467 & ~n21492 ;
  assign n21491 = n21467 ^ n21462 ;
  assign n21493 = n21492 ^ n21491 ;
  assign n21494 = x185 & ~n21493 ;
  assign n21496 = n21495 ^ n21494 ;
  assign n21483 = n21458 ^ n21157 ;
  assign n21484 = n21457 & ~n21483 ;
  assign n21480 = n21198 ^ n20415 ;
  assign n21481 = n21480 ^ n20416 ;
  assign n21482 = n21481 ^ n21458 ;
  assign n21485 = n21484 ^ n21482 ;
  assign n21486 = n21485 ^ n21198 ;
  assign n21487 = n21486 ^ n20442 ;
  assign n21488 = n21487 ^ n19277 ;
  assign n21479 = n19260 ^ x184 ;
  assign n21489 = n21488 ^ n21479 ;
  assign n21476 = n21461 ^ n21451 ;
  assign n21477 = n21461 ^ n19260 ;
  assign n21478 = ~n21476 & n21477 ;
  assign n21490 = n21489 ^ n21478 ;
  assign n21497 = n21496 ^ n21490 ;
  assign n21474 = n20598 ^ n20581 ;
  assign n21498 = n21497 ^ n21474 ;
  assign n21475 = n21474 ^ n21445 ;
  assign n21499 = n21498 ^ n21475 ;
  assign n21500 = n21473 & ~n21499 ;
  assign n21501 = n21500 ^ n21475 ;
  assign n21503 = n20636 ^ n20600 ;
  assign n21504 = n21503 ^ n20621 ;
  assign n21506 = n21504 ^ n21474 ;
  assign n21502 = n20419 ^ x167 ;
  assign n21505 = n21504 ^ n21502 ;
  assign n21507 = n21506 ^ n21505 ;
  assign n21508 = ~n21501 & ~n21507 ;
  assign n21509 = n21508 ^ n21506 ;
  assign n21573 = n20682 ^ n20664 ;
  assign n21575 = n21573 ^ n20547 ;
  assign n21574 = n21573 ^ n21504 ;
  assign n21576 = n21575 ^ n21574 ;
  assign n21577 = ~n21509 & ~n21576 ;
  assign n21578 = n21577 ^ n21575 ;
  assign n21579 = n20548 ^ n20547 ;
  assign n21590 = n21579 ^ n21573 ;
  assign n21591 = ~n21578 & n21590 ;
  assign n21588 = n20725 ^ n20708 ;
  assign n21589 = n21588 ^ n21573 ;
  assign n21592 = n21591 ^ n21589 ;
  assign n21593 = n20549 ^ n20545 ;
  assign n21628 = n21593 ^ n21588 ;
  assign n21629 = ~n21592 & ~n21628 ;
  assign n21630 = n21629 ^ n21593 ;
  assign n21632 = n21631 ^ n21630 ;
  assign n21649 = n21630 ^ n21627 ;
  assign n21650 = ~n21632 & n21649 ;
  assign n21654 = n21653 ^ n21650 ;
  assign n21670 = n20851 ^ n20834 ;
  assign n21671 = n21670 ^ n21652 ;
  assign n21672 = n21671 ^ n21670 ;
  assign n21648 = n20630 ^ n20590 ;
  assign n21673 = n21672 ^ n21648 ;
  assign n21674 = n21654 & n21673 ;
  assign n21675 = n21674 ^ n21671 ;
  assign n21692 = n20892 ^ n20853 ;
  assign n21693 = n21692 ^ n20877 ;
  assign n21695 = n21693 ^ n21670 ;
  assign n21676 = n20673 ^ n20631 ;
  assign n21694 = n21693 ^ n21676 ;
  assign n21696 = n21695 ^ n21694 ;
  assign n21697 = ~n21675 & ~n21696 ;
  assign n21698 = n21697 ^ n21695 ;
  assign n21715 = n20939 ^ n20917 ;
  assign n21717 = n21715 ^ n21693 ;
  assign n21699 = n20717 ^ n20674 ;
  assign n21716 = n21715 ^ n21699 ;
  assign n21718 = n21717 ^ n21716 ;
  assign n21719 = ~n21698 & ~n21718 ;
  assign n21720 = n21719 ^ n21717 ;
  assign n21737 = n20974 ^ n20941 ;
  assign n21738 = n21737 ^ n20962 ;
  assign n21740 = n21738 ^ n21715 ;
  assign n21721 = n20759 ^ n20718 ;
  assign n21739 = n21738 ^ n21721 ;
  assign n21741 = n21740 ^ n21739 ;
  assign n21742 = n21720 & ~n21741 ;
  assign n21743 = n21742 ^ n21740 ;
  assign n21760 = n21018 ^ n21001 ;
  assign n21762 = n21760 ^ n21738 ;
  assign n21744 = n20801 ^ n20760 ;
  assign n21761 = n21760 ^ n21744 ;
  assign n21763 = n21762 ^ n21761 ;
  assign n21764 = ~n21743 & ~n21763 ;
  assign n21765 = n21764 ^ n21762 ;
  assign n21781 = n21045 ^ n20520 ;
  assign n21783 = n21781 ^ n21760 ;
  assign n21766 = n20843 ^ n20802 ;
  assign n21782 = n21781 ^ n21766 ;
  assign n21784 = n21783 ^ n21782 ;
  assign n21785 = n21765 & n21784 ;
  assign n21786 = n21785 ^ n21783 ;
  assign n21807 = n21099 ^ n21086 ;
  assign n21808 = n21807 ^ n21083 ;
  assign n21810 = n21808 ^ n21781 ;
  assign n21787 = n20886 ^ n20844 ;
  assign n21809 = n21808 ^ n21787 ;
  assign n21811 = n21810 ^ n21809 ;
  assign n21812 = n21786 & n21811 ;
  assign n21813 = n21812 ^ n21810 ;
  assign n21815 = n21814 ^ n21813 ;
  assign n21816 = n21815 ^ n21087 ;
  assign n21767 = n21766 ^ n21765 ;
  assign n21768 = n21767 ^ n21002 ;
  assign n21790 = n21768 ^ n19591 ;
  assign n21745 = n21744 ^ n21743 ;
  assign n21746 = n21745 ^ n20963 ;
  assign n21755 = n21746 ^ n19596 ;
  assign n21722 = n21721 ^ n21720 ;
  assign n21723 = n21722 ^ n20918 ;
  assign n21732 = n21723 ^ n20383 ;
  assign n21700 = n21699 ^ n21698 ;
  assign n21701 = n21700 ^ n20878 ;
  assign n21710 = n21701 ^ n19601 ;
  assign n21677 = n21676 ^ n21675 ;
  assign n21678 = n21677 ^ n20835 ;
  assign n21687 = n21678 ^ n19606 ;
  assign n21655 = n21654 ^ n21648 ;
  assign n21656 = n21655 ^ n20793 ;
  assign n21665 = n21656 ^ n19611 ;
  assign n21633 = n21632 ^ n21627 ;
  assign n21634 = n21633 ^ n20751 ;
  assign n21643 = n21634 ^ n20220 ;
  assign n21512 = n21502 ^ n21501 ;
  assign n21513 = n21512 ^ n20582 ;
  assign n21514 = n21513 ^ n20051 ;
  assign n21515 = n21497 ^ n21473 ;
  assign n21516 = n21515 ^ n20537 ;
  assign n21517 = n21516 ^ n20010 ;
  assign n21526 = n21469 ^ n21444 ;
  assign n21527 = n21526 ^ n20494 ;
  assign n21520 = n21439 ^ n21415 ;
  assign n21521 = n21520 ^ n20465 ;
  assign n21518 = n21411 ^ n19922 ;
  assign n21519 = n19923 & n21518 ;
  assign n21522 = n21521 ^ n21519 ;
  assign n21523 = n21521 ^ n19927 ;
  assign n21524 = n21522 & n21523 ;
  assign n21525 = n21524 ^ n19927 ;
  assign n21528 = n21527 ^ n21525 ;
  assign n21529 = n21527 ^ n19967 ;
  assign n21530 = ~n21528 & n21529 ;
  assign n21531 = n21530 ^ n19967 ;
  assign n21532 = n21531 ^ n21516 ;
  assign n21533 = n21517 & n21532 ;
  assign n21534 = n21533 ^ n20010 ;
  assign n21535 = n21534 ^ n21513 ;
  assign n21536 = ~n21514 & n21535 ;
  assign n21537 = n21536 ^ n20051 ;
  assign n21538 = n21537 ^ n20094 ;
  assign n21510 = n21509 ^ n20547 ;
  assign n21511 = n21510 ^ n20622 ;
  assign n21582 = n21537 ^ n21511 ;
  assign n21583 = ~n21538 & n21582 ;
  assign n21584 = n21583 ^ n20094 ;
  assign n21585 = n21584 ^ n20138 ;
  assign n21580 = n21579 ^ n21578 ;
  assign n21581 = n21580 ^ n20665 ;
  assign n21596 = n21584 ^ n21581 ;
  assign n21597 = ~n21585 & ~n21596 ;
  assign n21598 = n21597 ^ n20138 ;
  assign n21599 = n21598 ^ n20177 ;
  assign n21594 = n21593 ^ n21592 ;
  assign n21595 = n21594 ^ n20709 ;
  assign n21622 = n21598 ^ n21595 ;
  assign n21623 = n21599 & ~n21622 ;
  assign n21624 = n21623 ^ n20177 ;
  assign n21644 = n21634 ^ n21624 ;
  assign n21645 = ~n21643 & ~n21644 ;
  assign n21646 = n21645 ^ n20220 ;
  assign n21666 = n21656 ^ n21646 ;
  assign n21667 = ~n21665 & n21666 ;
  assign n21668 = n21667 ^ n19611 ;
  assign n21688 = n21678 ^ n21668 ;
  assign n21689 = ~n21687 & ~n21688 ;
  assign n21690 = n21689 ^ n19606 ;
  assign n21711 = n21701 ^ n21690 ;
  assign n21712 = ~n21710 & ~n21711 ;
  assign n21713 = n21712 ^ n19601 ;
  assign n21733 = n21723 ^ n21713 ;
  assign n21734 = n21732 & ~n21733 ;
  assign n21735 = n21734 ^ n20383 ;
  assign n21756 = n21746 ^ n21735 ;
  assign n21757 = ~n21755 & n21756 ;
  assign n21758 = n21757 ^ n19596 ;
  assign n21791 = n21768 ^ n21758 ;
  assign n21792 = ~n21790 & ~n21791 ;
  assign n21793 = n21792 ^ n19591 ;
  assign n21794 = n21793 ^ n19697 ;
  assign n21788 = n21787 ^ n21786 ;
  assign n21789 = n21788 ^ n21045 ;
  assign n21803 = n21793 ^ n21789 ;
  assign n21804 = ~n21794 & n21803 ;
  assign n21805 = n21804 ^ n19697 ;
  assign n21806 = n21805 ^ n19811 ;
  assign n21817 = n21816 ^ n21806 ;
  assign n21795 = n21794 ^ n21789 ;
  assign n21798 = n21795 ^ x264 ;
  assign n21586 = n21585 ^ n21581 ;
  assign n21539 = n21538 ^ n21511 ;
  assign n21540 = n21539 ^ x258 ;
  assign n21543 = x263 & ~n21518 ;
  assign n21541 = n21519 ^ n19927 ;
  assign n21542 = n21541 ^ n21521 ;
  assign n21544 = n21543 ^ n21542 ;
  assign n21545 = n21525 ^ n19967 ;
  assign n21546 = n21545 ^ n21527 ;
  assign n21547 = n21546 ^ x262 ;
  assign n21548 = n21547 ^ n21542 ;
  assign n21549 = n21548 ^ n21546 ;
  assign n21550 = ~n21544 & n21549 ;
  assign n21551 = n21550 ^ n21547 ;
  assign n21552 = n21531 ^ n20010 ;
  assign n21553 = n21552 ^ n21516 ;
  assign n21555 = n21553 ^ x261 ;
  assign n21554 = n21553 ^ n21546 ;
  assign n21556 = n21555 ^ n21554 ;
  assign n21557 = n21551 & ~n21556 ;
  assign n21558 = n21557 ^ n21555 ;
  assign n21559 = n21534 ^ n20051 ;
  assign n21560 = n21559 ^ n21513 ;
  assign n21562 = n21560 ^ x260 ;
  assign n21561 = n21560 ^ n21553 ;
  assign n21563 = n21562 ^ n21561 ;
  assign n21564 = n21558 & ~n21563 ;
  assign n21565 = n21564 ^ n21562 ;
  assign n21567 = n21539 ^ x259 ;
  assign n21566 = n21560 ^ n21539 ;
  assign n21568 = n21567 ^ n21566 ;
  assign n21569 = n21565 & ~n21568 ;
  assign n21570 = n21569 ^ n21567 ;
  assign n21571 = n21540 & ~n21570 ;
  assign n21572 = n21571 ^ x258 ;
  assign n21587 = n21586 ^ n21572 ;
  assign n21600 = n21599 ^ n21595 ;
  assign n21601 = n21600 ^ x257 ;
  assign n21602 = n21601 ^ n21572 ;
  assign n21603 = n21602 ^ n21600 ;
  assign n21604 = ~n21587 & n21603 ;
  assign n21605 = n21604 ^ n21601 ;
  assign n21625 = n21624 ^ n20220 ;
  assign n21635 = n21634 ^ n21625 ;
  assign n21637 = n21635 ^ x256 ;
  assign n21636 = n21635 ^ n21600 ;
  assign n21638 = n21637 ^ n21636 ;
  assign n21639 = ~n21605 & n21638 ;
  assign n21640 = n21639 ^ n21637 ;
  assign n21647 = n21646 ^ n19611 ;
  assign n21657 = n21656 ^ n21647 ;
  assign n21659 = n21657 ^ x271 ;
  assign n21658 = n21657 ^ n21635 ;
  assign n21660 = n21659 ^ n21658 ;
  assign n21661 = n21640 & ~n21660 ;
  assign n21662 = n21661 ^ n21659 ;
  assign n21669 = n21668 ^ n19606 ;
  assign n21679 = n21678 ^ n21669 ;
  assign n21681 = n21679 ^ x270 ;
  assign n21680 = n21679 ^ n21657 ;
  assign n21682 = n21681 ^ n21680 ;
  assign n21683 = ~n21662 & n21682 ;
  assign n21684 = n21683 ^ n21681 ;
  assign n21691 = n21690 ^ n19601 ;
  assign n21702 = n21701 ^ n21691 ;
  assign n21704 = n21702 ^ x269 ;
  assign n21703 = n21702 ^ n21679 ;
  assign n21705 = n21704 ^ n21703 ;
  assign n21706 = ~n21684 & n21705 ;
  assign n21707 = n21706 ^ n21704 ;
  assign n21714 = n21713 ^ n20383 ;
  assign n21724 = n21723 ^ n21714 ;
  assign n21726 = n21724 ^ x268 ;
  assign n21725 = n21724 ^ n21702 ;
  assign n21727 = n21726 ^ n21725 ;
  assign n21728 = n21707 & ~n21727 ;
  assign n21729 = n21728 ^ n21726 ;
  assign n21736 = n21735 ^ n19596 ;
  assign n21747 = n21746 ^ n21736 ;
  assign n21749 = n21747 ^ x267 ;
  assign n21748 = n21747 ^ n21724 ;
  assign n21750 = n21749 ^ n21748 ;
  assign n21751 = n21729 & ~n21750 ;
  assign n21752 = n21751 ^ n21749 ;
  assign n21759 = n21758 ^ n19591 ;
  assign n21769 = n21768 ^ n21759 ;
  assign n21771 = n21769 ^ x266 ;
  assign n21770 = n21769 ^ n21747 ;
  assign n21772 = n21771 ^ n21770 ;
  assign n21773 = ~n21752 & n21772 ;
  assign n21774 = n21773 ^ n21771 ;
  assign n21777 = n21769 ^ x265 ;
  assign n21778 = ~n21774 & n21777 ;
  assign n21779 = n21778 ^ x265 ;
  assign n21799 = n21795 ^ n21779 ;
  assign n21800 = n21798 & ~n21799 ;
  assign n21801 = n21800 ^ x264 ;
  assign n21820 = n21817 ^ n21801 ;
  assign n21821 = n21816 ^ n21805 ;
  assign n21828 = n20966 ^ n20927 ;
  assign n21822 = n21171 ^ n21129 ;
  assign n21824 = n21822 ^ n21808 ;
  assign n21823 = n21822 ^ n21814 ;
  assign n21825 = n21824 ^ n21823 ;
  assign n21826 = n21813 & n21825 ;
  assign n21827 = n21826 ^ n21824 ;
  assign n21829 = n21828 ^ n21827 ;
  assign n21830 = n21829 ^ n21129 ;
  assign n21831 = n21830 ^ n19811 ;
  assign n21832 = n21831 ^ n21805 ;
  assign n21833 = n21832 ^ n21830 ;
  assign n21834 = n21821 & ~n21833 ;
  assign n21835 = n21834 ^ n21831 ;
  assign n21836 = n21835 ^ n20646 ;
  assign n21837 = n21836 ^ x279 ;
  assign n21838 = n21837 ^ n21801 ;
  assign n21839 = n21838 ^ n21836 ;
  assign n21840 = n21820 & n21839 ;
  assign n21841 = n21840 ^ n21837 ;
  assign n21850 = n21010 ^ n20967 ;
  assign n21844 = n21174 ^ n20653 ;
  assign n21846 = n21844 ^ n21822 ;
  assign n21845 = n21844 ^ n21828 ;
  assign n21847 = n21846 ^ n21845 ;
  assign n21848 = n21827 & n21847 ;
  assign n21849 = n21848 ^ n21846 ;
  assign n21851 = n21850 ^ n21849 ;
  assign n21852 = n21851 ^ n21174 ;
  assign n21854 = n21852 ^ n20646 ;
  assign n21853 = n21852 ^ n21830 ;
  assign n21855 = n21854 ^ n21853 ;
  assign n21856 = n21835 & n21855 ;
  assign n21857 = n21856 ^ n21854 ;
  assign n21858 = n21857 ^ n19846 ;
  assign n21860 = n21858 ^ x278 ;
  assign n21859 = n21858 ^ n21836 ;
  assign n21861 = n21860 ^ n21859 ;
  assign n21862 = ~n21841 & n21861 ;
  assign n21863 = n21862 ^ n21860 ;
  assign n21875 = n21852 ^ n19846 ;
  assign n21876 = n21857 & n21875 ;
  assign n21877 = n21876 ^ n19846 ;
  assign n21878 = n21877 ^ n19870 ;
  assign n21872 = n21053 ^ n21011 ;
  assign n21866 = n21229 ^ n21207 ;
  assign n21868 = n21866 ^ n21844 ;
  assign n21867 = n21866 ^ n21850 ;
  assign n21869 = n21868 ^ n21867 ;
  assign n21870 = n21849 & n21869 ;
  assign n21871 = n21870 ^ n21868 ;
  assign n21873 = n21872 ^ n21871 ;
  assign n21874 = n21873 ^ n21211 ;
  assign n21879 = n21878 ^ n21874 ;
  assign n21881 = n21879 ^ x277 ;
  assign n21880 = n21879 ^ n21858 ;
  assign n21882 = n21881 ^ n21880 ;
  assign n21883 = n21863 & ~n21882 ;
  assign n21884 = n21883 ^ n21881 ;
  assign n21896 = n21877 ^ n21874 ;
  assign n21897 = ~n21878 & ~n21896 ;
  assign n21898 = n21897 ^ n19870 ;
  assign n21899 = n21898 ^ n19951 ;
  assign n21893 = n21095 ^ n21054 ;
  assign n21887 = n21233 ^ n20738 ;
  assign n21889 = n21887 ^ n21866 ;
  assign n21888 = n21887 ^ n21872 ;
  assign n21890 = n21889 ^ n21888 ;
  assign n21891 = ~n21871 & n21890 ;
  assign n21892 = n21891 ^ n21889 ;
  assign n21894 = n21893 ^ n21892 ;
  assign n21895 = n21894 ^ n21233 ;
  assign n21900 = n21899 ^ n21895 ;
  assign n21902 = n21900 ^ x276 ;
  assign n21901 = n21900 ^ n21879 ;
  assign n21903 = n21902 ^ n21901 ;
  assign n21904 = n21884 & ~n21903 ;
  assign n21905 = n21904 ^ n21902 ;
  assign n21917 = n21898 ^ n21895 ;
  assign n21918 = ~n21899 & ~n21917 ;
  assign n21919 = n21918 ^ n19951 ;
  assign n21920 = n21919 ^ n19994 ;
  assign n21914 = n21142 ^ n21096 ;
  assign n21910 = n20780 ^ n20397 ;
  assign n21911 = n21910 ^ n21250 ;
  assign n21912 = n21911 ^ n21887 ;
  assign n21908 = n21893 ^ n21887 ;
  assign n21909 = ~n21892 & n21908 ;
  assign n21913 = n21912 ^ n21909 ;
  assign n21915 = n21914 ^ n21913 ;
  assign n21916 = n21915 ^ n21251 ;
  assign n21921 = n21920 ^ n21916 ;
  assign n21923 = n21921 ^ x275 ;
  assign n21922 = n21921 ^ n21900 ;
  assign n21924 = n21923 ^ n21922 ;
  assign n21925 = ~n21905 & n21924 ;
  assign n21926 = n21925 ^ n21923 ;
  assign n21927 = n21926 ^ x274 ;
  assign n21606 = n21605 ^ x256 ;
  assign n21607 = n21551 ^ x261 ;
  assign n21608 = n21518 ^ x263 ;
  assign n21609 = n21543 ^ x262 ;
  assign n21610 = n21609 ^ n21542 ;
  assign n21611 = ~n21608 & n21610 ;
  assign n21612 = ~n21607 & n21611 ;
  assign n21613 = n21558 ^ x260 ;
  assign n21614 = n21612 & ~n21613 ;
  assign n21615 = n21565 ^ x259 ;
  assign n21616 = n21614 & ~n21615 ;
  assign n21617 = n21570 ^ x258 ;
  assign n21618 = n21616 & n21617 ;
  assign n21619 = n21587 ^ x257 ;
  assign n21620 = n21618 & n21619 ;
  assign n21621 = ~n21606 & ~n21620 ;
  assign n21641 = n21640 ^ x271 ;
  assign n21642 = ~n21621 & ~n21641 ;
  assign n21663 = n21662 ^ x270 ;
  assign n21664 = ~n21642 & ~n21663 ;
  assign n21685 = n21684 ^ x269 ;
  assign n21686 = n21664 & ~n21685 ;
  assign n21708 = n21707 ^ x268 ;
  assign n21709 = ~n21686 & ~n21708 ;
  assign n21730 = n21729 ^ x267 ;
  assign n21731 = ~n21709 & n21730 ;
  assign n21753 = n21752 ^ x266 ;
  assign n21754 = n21731 & ~n21753 ;
  assign n21775 = n21774 ^ x265 ;
  assign n21776 = n21754 & ~n21775 ;
  assign n21780 = n21779 ^ x264 ;
  assign n21796 = n21795 ^ n21780 ;
  assign n21797 = n21776 & ~n21796 ;
  assign n21802 = n21801 ^ x279 ;
  assign n21818 = n21817 ^ n21802 ;
  assign n21819 = n21797 & n21818 ;
  assign n21842 = n21841 ^ x278 ;
  assign n21843 = ~n21819 & n21842 ;
  assign n21864 = n21863 ^ x277 ;
  assign n21865 = n21843 & ~n21864 ;
  assign n21885 = n21884 ^ x276 ;
  assign n21886 = n21865 & ~n21885 ;
  assign n21906 = n21905 ^ x275 ;
  assign n21907 = ~n21886 & ~n21906 ;
  assign n21928 = n21927 ^ n21907 ;
  assign n21955 = n21928 ^ n20418 ;
  assign n21956 = n20463 & n21955 ;
  assign n21929 = n21412 ^ n21411 ;
  assign n21952 = ~n21928 & ~n21929 ;
  assign n21940 = n21919 ^ n21916 ;
  assign n21941 = ~n21920 & ~n21940 ;
  assign n21942 = n21941 ^ n19994 ;
  assign n21943 = n21942 ^ n20036 ;
  assign n21932 = n21184 ^ n21143 ;
  assign n21933 = n21932 ^ n21914 ;
  assign n21934 = n21933 ^ n21911 ;
  assign n21935 = n21934 ^ n21932 ;
  assign n21936 = ~n21913 & ~n21935 ;
  assign n21937 = n21936 ^ n21933 ;
  assign n21938 = n21937 ^ n21273 ;
  assign n21939 = n21938 ^ n21274 ;
  assign n21944 = n21943 ^ n21939 ;
  assign n21946 = n21944 ^ x274 ;
  assign n21945 = n21944 ^ n21921 ;
  assign n21947 = n21946 ^ n21945 ;
  assign n21948 = n21926 & ~n21947 ;
  assign n21949 = n21948 ^ n21946 ;
  assign n21950 = n21949 ^ x273 ;
  assign n21931 = n21907 & n21927 ;
  assign n21951 = n21950 ^ n21931 ;
  assign n21953 = n21952 ^ n21951 ;
  assign n21954 = n21953 ^ n21414 ;
  assign n21957 = n21956 ^ n21954 ;
  assign n21989 = n21956 ^ n20471 ;
  assign n21990 = n21957 & ~n21989 ;
  assign n21991 = n21990 ^ n20471 ;
  assign n21992 = n21991 ^ n20510 ;
  assign n21984 = n21952 ^ n21520 ;
  assign n21985 = ~n21953 & ~n21984 ;
  assign n21986 = n21985 ^ n21520 ;
  assign n21978 = n21944 ^ x273 ;
  assign n21979 = ~n21949 & n21978 ;
  assign n21980 = n21979 ^ x273 ;
  assign n21981 = n21980 ^ x272 ;
  assign n21973 = n21942 ^ n21939 ;
  assign n21974 = ~n21943 & ~n21973 ;
  assign n21975 = n21974 ^ n20036 ;
  assign n21976 = n21975 ^ n20073 ;
  assign n21969 = n21294 ^ n21273 ;
  assign n21967 = n21932 ^ n21273 ;
  assign n21968 = n21937 & n21967 ;
  assign n21970 = n21969 ^ n21968 ;
  assign n21966 = n21223 ^ n21185 ;
  assign n21971 = n21970 ^ n21966 ;
  assign n21972 = n21971 ^ n21295 ;
  assign n21977 = n21976 ^ n21972 ;
  assign n21982 = n21981 ^ n21977 ;
  assign n21965 = n21931 & ~n21950 ;
  assign n21983 = n21982 ^ n21965 ;
  assign n21987 = n21986 ^ n21983 ;
  assign n21988 = n21987 ^ n21416 ;
  assign n21993 = n21992 ^ n21988 ;
  assign n21959 = x359 & ~n21955 ;
  assign n21958 = n21957 ^ n20471 ;
  assign n21960 = n21959 ^ n21958 ;
  assign n21962 = n21959 ^ x358 ;
  assign n21963 = ~n21960 & n21962 ;
  assign n21964 = n21963 ^ x358 ;
  assign n21994 = n21993 ^ n21964 ;
  assign n22022 = n21991 ^ n21988 ;
  assign n22023 = ~n21992 & ~n22022 ;
  assign n22024 = n22023 ^ n20510 ;
  assign n22025 = n22024 ^ n20556 ;
  assign n22014 = n21241 ^ n21224 ;
  assign n22009 = n21316 ^ n21294 ;
  assign n22010 = n22009 ^ n21316 ;
  assign n22011 = n22010 ^ n21966 ;
  assign n22012 = ~n21970 & ~n22011 ;
  assign n22013 = n22012 ^ n22009 ;
  assign n22015 = n22014 ^ n22013 ;
  assign n22016 = n22015 ^ n21317 ;
  assign n22005 = n21975 ^ n21972 ;
  assign n22006 = ~n21976 & ~n22005 ;
  assign n22007 = n22006 ^ n20073 ;
  assign n22008 = n22007 ^ n20122 ;
  assign n22017 = n22016 ^ n22008 ;
  assign n22001 = n21980 ^ n21977 ;
  assign n22002 = n21981 & n22001 ;
  assign n22003 = n22002 ^ x272 ;
  assign n22004 = n22003 ^ x287 ;
  assign n22018 = n22017 ^ n22004 ;
  assign n22000 = ~n21965 & ~n21982 ;
  assign n22019 = n22018 ^ n22000 ;
  assign n21997 = n21986 ^ n21526 ;
  assign n21998 = n21987 & n21997 ;
  assign n21999 = n21998 ^ n21526 ;
  assign n22020 = n22019 ^ n21999 ;
  assign n22021 = n22020 ^ n21445 ;
  assign n22026 = n22025 ^ n22021 ;
  assign n22028 = n22026 ^ x357 ;
  assign n22027 = n22026 ^ n21964 ;
  assign n22029 = n22028 ^ n22027 ;
  assign n22030 = ~n21994 & n22029 ;
  assign n22031 = n22030 ^ n22028 ;
  assign n22069 = n22026 ^ x356 ;
  assign n22070 = ~n22031 & n22069 ;
  assign n22071 = n22070 ^ x356 ;
  assign n22064 = n22024 ^ n22021 ;
  assign n22065 = ~n22025 & n22064 ;
  assign n22066 = n22065 ^ n20556 ;
  assign n22067 = n22066 ^ n20596 ;
  assign n22038 = n22017 ^ n22003 ;
  assign n22039 = n22016 ^ n22007 ;
  assign n22046 = n21259 ^ n21242 ;
  assign n22040 = n21348 ^ n21333 ;
  assign n22042 = n22040 ^ n21316 ;
  assign n22041 = n22040 ^ n22014 ;
  assign n22043 = n22042 ^ n22041 ;
  assign n22044 = ~n22013 & n22043 ;
  assign n22045 = n22044 ^ n22042 ;
  assign n22047 = n22046 ^ n22045 ;
  assign n22048 = n22047 ^ n21333 ;
  assign n22049 = n22048 ^ n20122 ;
  assign n22050 = n22049 ^ n22007 ;
  assign n22051 = n22050 ^ n22048 ;
  assign n22052 = ~n22039 & n22051 ;
  assign n22053 = n22052 ^ n22049 ;
  assign n22054 = n22053 ^ n20983 ;
  assign n22055 = n22054 ^ x287 ;
  assign n22056 = n22055 ^ n22003 ;
  assign n22057 = n22056 ^ n22054 ;
  assign n22058 = n22038 & n22057 ;
  assign n22059 = n22058 ^ n22055 ;
  assign n22060 = n22059 ^ x286 ;
  assign n22037 = ~n22000 & n22018 ;
  assign n22061 = n22060 ^ n22037 ;
  assign n22034 = n22019 ^ n21515 ;
  assign n22035 = n22020 & ~n22034 ;
  assign n22036 = n22035 ^ n21515 ;
  assign n22062 = n22061 ^ n22036 ;
  assign n22063 = n22062 ^ n21474 ;
  assign n22068 = n22067 ^ n22063 ;
  assign n22072 = n22071 ^ n22068 ;
  assign n22103 = n22066 ^ n22063 ;
  assign n22104 = n22067 & n22103 ;
  assign n22105 = n22104 ^ n20596 ;
  assign n22106 = n22105 ^ n20636 ;
  assign n22098 = n22061 ^ n21512 ;
  assign n22099 = n22062 & ~n22098 ;
  assign n22100 = n22099 ^ n21512 ;
  assign n22082 = n21281 ^ n21260 ;
  assign n22076 = n21355 ^ n20989 ;
  assign n22078 = n22076 ^ n22040 ;
  assign n22077 = n22076 ^ n22046 ;
  assign n22079 = n22078 ^ n22077 ;
  assign n22080 = ~n22045 & ~n22079 ;
  assign n22081 = n22080 ^ n22078 ;
  assign n22083 = n22082 ^ n22081 ;
  assign n22084 = n22083 ^ n21355 ;
  assign n22086 = n22084 ^ n20983 ;
  assign n22085 = n22084 ^ n22048 ;
  assign n22087 = n22086 ^ n22085 ;
  assign n22088 = n22053 & ~n22087 ;
  assign n22089 = n22088 ^ n22086 ;
  assign n22090 = n22089 ^ n20204 ;
  assign n22092 = n22090 ^ x286 ;
  assign n22091 = n22090 ^ n22054 ;
  assign n22093 = n22092 ^ n22091 ;
  assign n22094 = ~n22059 & n22093 ;
  assign n22095 = n22094 ^ n22092 ;
  assign n22096 = n22095 ^ x285 ;
  assign n22075 = n22037 & ~n22060 ;
  assign n22097 = n22096 ^ n22075 ;
  assign n22101 = n22100 ^ n22097 ;
  assign n22102 = n22101 ^ n21504 ;
  assign n22107 = n22106 ^ n22102 ;
  assign n22108 = n22107 ^ x355 ;
  assign n22109 = n22108 ^ n22071 ;
  assign n22110 = n22109 ^ n22107 ;
  assign n22111 = ~n22072 & n22110 ;
  assign n22112 = n22111 ^ n22108 ;
  assign n22140 = n22105 ^ n22102 ;
  assign n22141 = ~n22106 & ~n22140 ;
  assign n22142 = n22141 ^ n20636 ;
  assign n22143 = n22142 ^ n20680 ;
  assign n22125 = n22082 ^ n22076 ;
  assign n22126 = ~n22081 & ~n22125 ;
  assign n22124 = n22076 ^ n21379 ;
  assign n22127 = n22126 ^ n22124 ;
  assign n22123 = n21303 ^ n21282 ;
  assign n22128 = n22127 ^ n22123 ;
  assign n22129 = n22128 ^ n21380 ;
  assign n22119 = n22084 ^ n20204 ;
  assign n22120 = n22089 & n22119 ;
  assign n22121 = n22120 ^ n20204 ;
  assign n22122 = n22121 ^ n20246 ;
  assign n22130 = n22129 ^ n22122 ;
  assign n22132 = n22130 ^ x285 ;
  assign n22131 = n22130 ^ n22090 ;
  assign n22133 = n22132 ^ n22131 ;
  assign n22134 = n22095 & ~n22133 ;
  assign n22135 = n22134 ^ n22132 ;
  assign n22136 = n22135 ^ x284 ;
  assign n22118 = n22075 & n22096 ;
  assign n22137 = n22136 ^ n22118 ;
  assign n22115 = n22100 ^ n21510 ;
  assign n22116 = ~n22101 & ~n22115 ;
  assign n22117 = n22116 ^ n21510 ;
  assign n22138 = n22137 ^ n22117 ;
  assign n22139 = n22138 ^ n21573 ;
  assign n22144 = n22143 ^ n22139 ;
  assign n22146 = n22144 ^ x354 ;
  assign n22145 = n22144 ^ n22107 ;
  assign n22147 = n22146 ^ n22145 ;
  assign n22148 = ~n22112 & n22147 ;
  assign n22149 = n22148 ^ n22146 ;
  assign n22179 = n22142 ^ n22139 ;
  assign n22180 = n22143 & n22179 ;
  assign n22181 = n22180 ^ n20680 ;
  assign n22182 = n22181 ^ n20723 ;
  assign n22175 = ~n22118 & ~n22136 ;
  assign n22165 = n21325 ^ n21304 ;
  assign n22160 = n21401 ^ n21379 ;
  assign n22161 = n22160 ^ n21401 ;
  assign n22162 = n22161 ^ n22123 ;
  assign n22163 = n22127 & ~n22162 ;
  assign n22164 = n22163 ^ n22160 ;
  assign n22166 = n22165 ^ n22164 ;
  assign n22167 = n22166 ^ n21402 ;
  assign n22155 = n22129 ^ n22121 ;
  assign n22156 = n22129 ^ n20246 ;
  assign n22157 = ~n22155 & ~n22156 ;
  assign n22158 = n22157 ^ n20246 ;
  assign n22159 = n22158 ^ n20285 ;
  assign n22168 = n22167 ^ n22159 ;
  assign n22170 = n22168 ^ x284 ;
  assign n22169 = n22168 ^ n22130 ;
  assign n22171 = n22170 ^ n22169 ;
  assign n22172 = n22135 & ~n22171 ;
  assign n22173 = n22172 ^ n22170 ;
  assign n22174 = n22173 ^ x283 ;
  assign n22176 = n22175 ^ n22174 ;
  assign n22152 = n22137 ^ n21580 ;
  assign n22153 = ~n22138 & n22152 ;
  assign n22154 = n22153 ^ n21580 ;
  assign n22177 = n22176 ^ n22154 ;
  assign n22178 = n22177 ^ n21588 ;
  assign n22183 = n22182 ^ n22178 ;
  assign n22185 = n22183 ^ x353 ;
  assign n22184 = n22183 ^ n22144 ;
  assign n22186 = n22185 ^ n22184 ;
  assign n22187 = n22149 & ~n22186 ;
  assign n22188 = n22187 ^ n22185 ;
  assign n22189 = n22188 ^ x352 ;
  assign n21961 = n21960 ^ x358 ;
  assign n21995 = n21994 ^ x357 ;
  assign n21996 = n21961 & n21995 ;
  assign n22032 = n22031 ^ x356 ;
  assign n22033 = n21996 & n22032 ;
  assign n22073 = n22072 ^ x355 ;
  assign n22074 = n22033 & n22073 ;
  assign n22113 = n22112 ^ x354 ;
  assign n22114 = ~n22074 & ~n22113 ;
  assign n22150 = n22149 ^ x353 ;
  assign n22151 = ~n22114 & ~n22150 ;
  assign n23238 = n22189 ^ n22151 ;
  assign n22204 = n21346 ^ n21326 ;
  assign n22200 = n21429 ^ n21401 ;
  assign n22199 = n22165 ^ n21429 ;
  assign n22201 = n22200 ^ n22199 ;
  assign n22202 = n22164 & n22201 ;
  assign n22203 = n22202 ^ n22200 ;
  assign n22205 = n22204 ^ n22203 ;
  assign n22206 = n22205 ^ n21430 ;
  assign n22194 = n22167 ^ n22158 ;
  assign n22195 = n22167 ^ n20285 ;
  assign n22196 = n22194 & n22195 ;
  assign n22197 = n22196 ^ n20285 ;
  assign n22198 = n22197 ^ n20327 ;
  assign n22207 = n22206 ^ n22198 ;
  assign n22209 = n22207 ^ x283 ;
  assign n22208 = n22207 ^ n22168 ;
  assign n22210 = n22209 ^ n22208 ;
  assign n22211 = n22173 & ~n22210 ;
  assign n22212 = n22211 ^ n22209 ;
  assign n22240 = n21367 ^ n21347 ;
  assign n22236 = n21459 ^ n21429 ;
  assign n22235 = n22204 ^ n21459 ;
  assign n22237 = n22236 ^ n22235 ;
  assign n22238 = n22203 & n22237 ;
  assign n22239 = n22238 ^ n22236 ;
  assign n22241 = n22240 ^ n22239 ;
  assign n22242 = n22241 ^ n21460 ;
  assign n22230 = n22206 ^ n22197 ;
  assign n22231 = n22206 ^ n20327 ;
  assign n22232 = n22230 & n22231 ;
  assign n22233 = n22232 ^ n20327 ;
  assign n22234 = n22233 ^ n20367 ;
  assign n22243 = n22242 ^ n22234 ;
  assign n22245 = n22243 ^ x282 ;
  assign n22244 = n22243 ^ n22207 ;
  assign n22246 = n22245 ^ n22244 ;
  assign n22247 = ~n22212 & n22246 ;
  assign n22248 = n22247 ^ n22245 ;
  assign n22213 = n22212 ^ x282 ;
  assign n22214 = ~n22174 & n22175 ;
  assign n22250 = n22213 & n22214 ;
  assign n22287 = n22250 ^ n22243 ;
  assign n22288 = ~n22248 & ~n22287 ;
  assign n22285 = n22250 ^ n22248 ;
  assign n22286 = ~x281 & n22285 ;
  assign n22289 = n22288 ^ n22286 ;
  assign n22279 = n22240 ^ n21459 ;
  assign n22280 = n22239 & ~n22279 ;
  assign n22276 = n21388 ^ n21368 ;
  assign n22277 = n22276 ^ n21485 ;
  assign n22278 = n22277 ^ n22240 ;
  assign n22281 = n22280 ^ n22278 ;
  assign n22282 = n22281 ^ n21487 ;
  assign n22275 = n20367 ^ x280 ;
  assign n22283 = n22282 ^ n22275 ;
  assign n22272 = n22242 ^ n22233 ;
  assign n22273 = n22242 ^ n20367 ;
  assign n22274 = n22272 & ~n22273 ;
  assign n22284 = n22283 ^ n22274 ;
  assign n22290 = n22289 ^ n22284 ;
  assign n22215 = n22214 ^ n22213 ;
  assign n22191 = n22176 ^ n21594 ;
  assign n22192 = n22177 & ~n22191 ;
  assign n22193 = n22192 ^ n21594 ;
  assign n22216 = n22215 ^ n22193 ;
  assign n22252 = n22215 ^ n21633 ;
  assign n22253 = ~n22216 & n22252 ;
  assign n22254 = n22253 ^ n21633 ;
  assign n22249 = n22248 ^ x281 ;
  assign n22251 = n22250 ^ n22249 ;
  assign n22255 = n22254 ^ n22251 ;
  assign n22269 = n22254 ^ n21655 ;
  assign n22270 = ~n22255 & n22269 ;
  assign n22271 = n22270 ^ n21655 ;
  assign n22291 = n22290 ^ n22271 ;
  assign n22309 = n22290 ^ n21677 ;
  assign n22310 = ~n22291 & ~n22309 ;
  assign n22311 = n22310 ^ n21677 ;
  assign n22327 = n22311 ^ n21700 ;
  assign n22328 = n21722 ^ n21608 ;
  assign n22329 = n22328 ^ n21722 ;
  assign n22330 = n22329 ^ n22311 ;
  assign n22331 = n22327 & ~n22330 ;
  assign n22332 = n22331 ^ n22328 ;
  assign n22333 = n21610 ^ n21608 ;
  assign n22350 = n22333 ^ n21722 ;
  assign n22351 = ~n22332 & n22350 ;
  assign n22349 = n21745 ^ n21722 ;
  assign n22352 = n22351 ^ n22349 ;
  assign n22370 = n21613 ^ n21612 ;
  assign n22353 = n21611 ^ n21607 ;
  assign n22371 = n22370 ^ n22353 ;
  assign n22372 = n22371 ^ n21745 ;
  assign n22373 = n22372 ^ n22370 ;
  assign n22374 = ~n22352 & n22373 ;
  assign n22375 = n22374 ^ n22371 ;
  assign n22386 = n21788 ^ n21767 ;
  assign n22385 = n22370 ^ n21788 ;
  assign n22387 = n22386 ^ n22385 ;
  assign n22388 = ~n22375 & n22387 ;
  assign n22389 = n22388 ^ n22386 ;
  assign n22390 = n21615 ^ n21614 ;
  assign n22410 = n22390 ^ n21788 ;
  assign n22411 = n22389 & n22410 ;
  assign n22412 = n22411 ^ n21788 ;
  assign n22408 = n21617 ^ n21616 ;
  assign n22437 = n22412 ^ n22408 ;
  assign n22438 = n21619 ^ n21618 ;
  assign n22439 = n22438 ^ n21815 ;
  assign n22440 = n22439 ^ n22408 ;
  assign n22441 = n22440 ^ n22438 ;
  assign n22442 = n22437 & ~n22441 ;
  assign n22443 = n22442 ^ n22439 ;
  assign n23120 = n22443 ^ n21829 ;
  assign n22218 = n22181 ^ n22178 ;
  assign n22219 = ~n22182 & ~n22218 ;
  assign n22220 = n22219 ^ n20723 ;
  assign n22221 = n22220 ^ n20766 ;
  assign n22217 = n22216 ^ n21627 ;
  assign n22222 = n22221 ^ n22217 ;
  assign n22224 = n22222 ^ x352 ;
  assign n22223 = n22222 ^ n22183 ;
  assign n22225 = n22224 ^ n22223 ;
  assign n22226 = n22188 & ~n22225 ;
  assign n22227 = n22226 ^ n22224 ;
  assign n22257 = n22220 ^ n22217 ;
  assign n22258 = ~n22221 & n22257 ;
  assign n22259 = n22258 ^ n20766 ;
  assign n22260 = n22259 ^ n20808 ;
  assign n22256 = n22255 ^ n21652 ;
  assign n22261 = n22260 ^ n22256 ;
  assign n22263 = n22261 ^ x367 ;
  assign n22262 = n22261 ^ n22222 ;
  assign n22264 = n22263 ^ n22262 ;
  assign n22265 = n22227 & ~n22264 ;
  assign n22266 = n22265 ^ n22263 ;
  assign n22293 = n22259 ^ n22256 ;
  assign n22294 = n22260 & ~n22293 ;
  assign n22295 = n22294 ^ n20808 ;
  assign n22296 = n22295 ^ n20849 ;
  assign n22292 = n22291 ^ n21670 ;
  assign n22297 = n22296 ^ n22292 ;
  assign n22299 = n22297 ^ x366 ;
  assign n22298 = n22297 ^ n22261 ;
  assign n22300 = n22299 ^ n22298 ;
  assign n22301 = ~n22266 & n22300 ;
  assign n22302 = n22301 ^ n22299 ;
  assign n22312 = n22311 ^ n21608 ;
  assign n22313 = n22312 ^ n21693 ;
  assign n22305 = n22295 ^ n22292 ;
  assign n22306 = ~n22296 & n22305 ;
  assign n22307 = n22306 ^ n20849 ;
  assign n22308 = n22307 ^ n20892 ;
  assign n22314 = n22313 ^ n22308 ;
  assign n22316 = n22314 ^ x365 ;
  assign n22315 = n22314 ^ n22297 ;
  assign n22317 = n22316 ^ n22315 ;
  assign n22318 = ~n22302 & n22317 ;
  assign n22319 = n22318 ^ n22316 ;
  assign n22338 = n22314 ^ x364 ;
  assign n22339 = ~n22319 & n22338 ;
  assign n22340 = n22339 ^ x364 ;
  assign n22334 = n22333 ^ n22332 ;
  assign n22335 = n22334 ^ n21722 ;
  assign n22336 = n22335 ^ n21715 ;
  assign n22322 = n22313 ^ n22307 ;
  assign n22323 = n22313 ^ n20892 ;
  assign n22324 = ~n22322 & ~n22323 ;
  assign n22325 = n22324 ^ n20892 ;
  assign n22326 = n22325 ^ n20937 ;
  assign n22337 = n22336 ^ n22326 ;
  assign n22341 = n22340 ^ n22337 ;
  assign n22354 = n22353 ^ n22352 ;
  assign n22355 = n22354 ^ n21745 ;
  assign n22356 = n22355 ^ n21738 ;
  assign n22344 = n22336 ^ n20937 ;
  assign n22345 = n22336 ^ n22325 ;
  assign n22346 = ~n22344 & n22345 ;
  assign n22347 = n22346 ^ n20937 ;
  assign n22348 = n22347 ^ n20974 ;
  assign n22357 = n22356 ^ n22348 ;
  assign n22358 = n22357 ^ x363 ;
  assign n22359 = n22358 ^ n22340 ;
  assign n22360 = n22359 ^ n22357 ;
  assign n22361 = n22341 & n22360 ;
  assign n22362 = n22361 ^ n22358 ;
  assign n22376 = n22375 ^ n21760 ;
  assign n22365 = n22356 ^ n20974 ;
  assign n22366 = n22356 ^ n22347 ;
  assign n22367 = ~n22365 & n22366 ;
  assign n22368 = n22367 ^ n20974 ;
  assign n22369 = n22368 ^ n21016 ;
  assign n22377 = n22376 ^ n22369 ;
  assign n22379 = n22377 ^ x362 ;
  assign n22378 = n22377 ^ n22357 ;
  assign n22380 = n22379 ^ n22378 ;
  assign n22381 = n22362 & ~n22380 ;
  assign n22382 = n22381 ^ n22379 ;
  assign n22394 = n22376 ^ n21016 ;
  assign n22395 = n22376 ^ n22368 ;
  assign n22396 = n22394 & n22395 ;
  assign n22397 = n22396 ^ n21016 ;
  assign n22398 = n22397 ^ n20520 ;
  assign n22391 = n22390 ^ n22389 ;
  assign n22392 = n22391 ^ n21788 ;
  assign n22393 = n22392 ^ n21781 ;
  assign n22399 = n22398 ^ n22393 ;
  assign n22401 = n22399 ^ x361 ;
  assign n22400 = n22399 ^ n22377 ;
  assign n22402 = n22401 ^ n22400 ;
  assign n22403 = ~n22382 & n22402 ;
  assign n22404 = n22403 ^ n22401 ;
  assign n22422 = n22399 ^ x360 ;
  assign n22423 = n22404 & ~n22422 ;
  assign n22424 = n22423 ^ x360 ;
  assign n22407 = n22397 ^ n22393 ;
  assign n22409 = n22408 ^ n21815 ;
  assign n22413 = n22412 ^ n22409 ;
  assign n22414 = n22413 ^ n21815 ;
  assign n22415 = n22414 ^ n21808 ;
  assign n22416 = n22415 ^ n20520 ;
  assign n22417 = n22416 ^ n22393 ;
  assign n22418 = n22417 ^ n22415 ;
  assign n22419 = ~n22407 & n22418 ;
  assign n22420 = n22419 ^ n22416 ;
  assign n22421 = n22420 ^ n21099 ;
  assign n22435 = n22424 ^ n22421 ;
  assign n22444 = n21822 ^ n21099 ;
  assign n22445 = n22444 ^ n22443 ;
  assign n22436 = n22415 ^ n21822 ;
  assign n22446 = n22445 ^ n22436 ;
  assign n22447 = n22446 ^ n22443 ;
  assign n22448 = n22420 & n22447 ;
  assign n22449 = n22448 ^ n22445 ;
  assign n22450 = n22449 ^ n21171 ;
  assign n22451 = n22450 ^ x375 ;
  assign n22452 = n22451 ^ n22421 ;
  assign n22453 = n22452 ^ n22450 ;
  assign n22454 = n22435 & ~n22453 ;
  assign n22455 = n22454 ^ n22451 ;
  assign n22479 = n22438 ^ n21829 ;
  assign n22480 = n22443 & ~n22479 ;
  assign n22478 = n21851 ^ n21829 ;
  assign n22481 = n22480 ^ n22478 ;
  assign n22477 = n21620 ^ n21606 ;
  assign n22482 = n22481 ^ n22477 ;
  assign n22483 = n22482 ^ n21851 ;
  assign n22484 = n22483 ^ n21844 ;
  assign n22485 = n22484 ^ n21171 ;
  assign n22475 = n22443 ^ n21129 ;
  assign n22476 = ~n22449 & ~n22475 ;
  assign n22486 = n22485 ^ n22476 ;
  assign n22487 = n22486 ^ n20653 ;
  assign n22489 = n22487 ^ x374 ;
  assign n22488 = n22487 ^ n22450 ;
  assign n22490 = n22489 ^ n22488 ;
  assign n22491 = n22455 & ~n22490 ;
  assign n22492 = n22491 ^ n22489 ;
  assign n22517 = n22483 ^ n21174 ;
  assign n22518 = ~n22486 & ~n22517 ;
  assign n22519 = n22518 ^ n20653 ;
  assign n22520 = n22519 ^ n20697 ;
  assign n22512 = n22477 ^ n21851 ;
  assign n22513 = n22481 & n22512 ;
  assign n22514 = n22513 ^ n21851 ;
  assign n22511 = n21641 ^ n21621 ;
  assign n22515 = n22514 ^ n22511 ;
  assign n22516 = n22515 ^ n21866 ;
  assign n22521 = n22520 ^ n22516 ;
  assign n22523 = n22521 ^ x373 ;
  assign n22522 = n22521 ^ n22487 ;
  assign n22524 = n22523 ^ n22522 ;
  assign n22525 = ~n22492 & n22524 ;
  assign n22526 = n22525 ^ n22523 ;
  assign n22559 = n22519 ^ n22516 ;
  assign n22560 = ~n22520 & n22559 ;
  assign n22561 = n22560 ^ n20697 ;
  assign n22562 = n22561 ^ n20738 ;
  assign n22555 = n21663 ^ n21642 ;
  assign n22551 = n21894 ^ n21873 ;
  assign n22550 = n22514 ^ n21894 ;
  assign n22552 = n22551 ^ n22550 ;
  assign n22553 = n22515 & n22552 ;
  assign n22554 = n22553 ^ n22551 ;
  assign n22556 = n22555 ^ n22554 ;
  assign n22557 = n22556 ^ n21894 ;
  assign n22558 = n22557 ^ n21887 ;
  assign n22563 = n22562 ^ n22558 ;
  assign n22565 = n22563 ^ x372 ;
  assign n22564 = n22563 ^ n22521 ;
  assign n22566 = n22565 ^ n22564 ;
  assign n22567 = ~n22526 & n22566 ;
  assign n22568 = n22567 ^ n22565 ;
  assign n22600 = n22561 ^ n22558 ;
  assign n22601 = ~n22562 & ~n22600 ;
  assign n22602 = n22601 ^ n20738 ;
  assign n22603 = n22602 ^ n20780 ;
  assign n22596 = n21685 ^ n21664 ;
  assign n22592 = n21915 ^ n21894 ;
  assign n22591 = n22555 ^ n21915 ;
  assign n22593 = n22592 ^ n22591 ;
  assign n22594 = ~n22554 & ~n22593 ;
  assign n22595 = n22594 ^ n22592 ;
  assign n22597 = n22596 ^ n22595 ;
  assign n22598 = n22597 ^ n21915 ;
  assign n22599 = n22598 ^ n21911 ;
  assign n22604 = n22603 ^ n22599 ;
  assign n22606 = n22604 ^ x371 ;
  assign n22605 = n22604 ^ n22563 ;
  assign n22607 = n22606 ^ n22605 ;
  assign n22608 = ~n22568 & n22607 ;
  assign n22609 = n22608 ^ n22606 ;
  assign n22641 = n22602 ^ n22599 ;
  assign n22642 = ~n22603 & n22641 ;
  assign n22643 = n22642 ^ n20780 ;
  assign n22644 = n22643 ^ n20822 ;
  assign n22637 = n21708 ^ n21686 ;
  assign n22633 = n21938 ^ n21915 ;
  assign n22632 = n22596 ^ n21938 ;
  assign n22634 = n22633 ^ n22632 ;
  assign n22635 = n22595 & n22634 ;
  assign n22636 = n22635 ^ n22633 ;
  assign n22638 = n22637 ^ n22636 ;
  assign n22639 = n22638 ^ n21938 ;
  assign n22640 = n22639 ^ n21273 ;
  assign n22645 = n22644 ^ n22640 ;
  assign n22647 = n22645 ^ x370 ;
  assign n22646 = n22645 ^ n22604 ;
  assign n22648 = n22647 ^ n22646 ;
  assign n22649 = ~n22609 & n22648 ;
  assign n22650 = n22649 ^ n22647 ;
  assign n22682 = n21730 ^ n21709 ;
  assign n22678 = n21971 ^ n21938 ;
  assign n22677 = n22637 ^ n21971 ;
  assign n22679 = n22678 ^ n22677 ;
  assign n22680 = n22636 & n22679 ;
  assign n22681 = n22680 ^ n22678 ;
  assign n22683 = n22682 ^ n22681 ;
  assign n22684 = n22683 ^ n21971 ;
  assign n22685 = n22684 ^ n21294 ;
  assign n22673 = n22643 ^ n22640 ;
  assign n22674 = ~n22644 & ~n22673 ;
  assign n22675 = n22674 ^ n20822 ;
  assign n22676 = n22675 ^ n20860 ;
  assign n22686 = n22685 ^ n22676 ;
  assign n22688 = n22686 ^ x369 ;
  assign n22687 = n22686 ^ n22645 ;
  assign n22689 = n22688 ^ n22687 ;
  assign n22690 = ~n22650 & n22689 ;
  assign n22691 = n22690 ^ n22688 ;
  assign n22729 = n22686 ^ x368 ;
  assign n22730 = ~n22691 & n22729 ;
  assign n22731 = n22730 ^ x368 ;
  assign n22714 = n22685 ^ n22675 ;
  assign n22717 = n22682 ^ n21971 ;
  assign n22718 = n22681 & n22717 ;
  assign n22719 = n22718 ^ n21971 ;
  assign n22715 = n21753 ^ n21731 ;
  assign n22716 = n22715 ^ n22015 ;
  assign n22720 = n22719 ^ n22716 ;
  assign n22721 = n22720 ^ n22015 ;
  assign n22722 = n22721 ^ n21316 ;
  assign n22723 = n22722 ^ n20860 ;
  assign n22724 = n22723 ^ n22675 ;
  assign n22725 = n22724 ^ n22722 ;
  assign n22726 = ~n22714 & n22725 ;
  assign n22727 = n22726 ^ n22723 ;
  assign n22728 = n22727 ^ n21310 ;
  assign n22754 = n22731 ^ n22728 ;
  assign n22763 = n22040 ^ n21310 ;
  assign n22760 = n21775 ^ n21754 ;
  assign n22756 = n22719 ^ n22715 ;
  assign n22757 = n22719 ^ n22015 ;
  assign n22758 = ~n22756 & n22757 ;
  assign n22759 = n22758 ^ n22015 ;
  assign n22761 = n22760 ^ n22759 ;
  assign n22764 = n22763 ^ n22761 ;
  assign n22755 = n22722 ^ n22040 ;
  assign n22762 = n22761 ^ n22755 ;
  assign n22765 = n22764 ^ n22762 ;
  assign n22766 = n22727 & ~n22765 ;
  assign n22767 = n22766 ^ n22764 ;
  assign n22768 = n22767 ^ n21348 ;
  assign n22769 = n22768 ^ x383 ;
  assign n22770 = n22769 ^ n22728 ;
  assign n22771 = n22770 ^ n22768 ;
  assign n22772 = n22754 & ~n22771 ;
  assign n22773 = n22772 ^ n22769 ;
  assign n22806 = n22761 ^ n21333 ;
  assign n22807 = ~n22767 & n22806 ;
  assign n22801 = n21796 ^ n21776 ;
  assign n22796 = n22083 ^ n22047 ;
  assign n22797 = n22796 ^ n22083 ;
  assign n22798 = n22797 ^ n22759 ;
  assign n22799 = ~n22761 & n22798 ;
  assign n22800 = n22799 ^ n22796 ;
  assign n22802 = n22801 ^ n22800 ;
  assign n22803 = n22802 ^ n22083 ;
  assign n22804 = n22803 ^ n22076 ;
  assign n22805 = n22804 ^ n21348 ;
  assign n22808 = n22807 ^ n22805 ;
  assign n22809 = n22808 ^ n20989 ;
  assign n22811 = n22809 ^ x382 ;
  assign n22810 = n22809 ^ n22768 ;
  assign n22812 = n22811 ^ n22810 ;
  assign n22813 = ~n22773 & n22812 ;
  assign n22814 = n22813 ^ n22811 ;
  assign n22846 = n21818 ^ n21797 ;
  assign n22842 = n22128 ^ n22083 ;
  assign n22841 = n22801 ^ n22128 ;
  assign n22843 = n22842 ^ n22841 ;
  assign n22844 = ~n22800 & ~n22843 ;
  assign n22845 = n22844 ^ n22842 ;
  assign n22847 = n22846 ^ n22845 ;
  assign n22848 = n22847 ^ n22128 ;
  assign n22849 = n22848 ^ n21379 ;
  assign n22837 = n22803 ^ n21355 ;
  assign n22838 = n22808 & ~n22837 ;
  assign n22839 = n22838 ^ n20989 ;
  assign n22840 = n22839 ^ n21031 ;
  assign n22850 = n22849 ^ n22840 ;
  assign n22852 = n22850 ^ x381 ;
  assign n22851 = n22850 ^ n22809 ;
  assign n22853 = n22852 ^ n22851 ;
  assign n22854 = n22814 & ~n22853 ;
  assign n22855 = n22854 ^ n22852 ;
  assign n22881 = n21842 ^ n21819 ;
  assign n22877 = n22166 ^ n22128 ;
  assign n22876 = n22846 ^ n22166 ;
  assign n22878 = n22877 ^ n22876 ;
  assign n22879 = ~n22845 & ~n22878 ;
  assign n22880 = n22879 ^ n22877 ;
  assign n22882 = n22881 ^ n22880 ;
  assign n22883 = n22882 ^ n22166 ;
  assign n22884 = n22883 ^ n21401 ;
  assign n22871 = n22849 ^ n22839 ;
  assign n22872 = n22849 ^ n21031 ;
  assign n22873 = n22871 & n22872 ;
  assign n22874 = n22873 ^ n21031 ;
  assign n22875 = n22874 ^ n21071 ;
  assign n22885 = n22884 ^ n22875 ;
  assign n22887 = n22885 ^ x380 ;
  assign n22886 = n22885 ^ n22850 ;
  assign n22888 = n22887 ^ n22886 ;
  assign n22889 = ~n22855 & n22888 ;
  assign n22890 = n22889 ^ n22887 ;
  assign n22919 = n21864 ^ n21843 ;
  assign n22915 = n22205 ^ n22166 ;
  assign n22914 = n22881 ^ n22205 ;
  assign n22916 = n22915 ^ n22914 ;
  assign n22917 = ~n22880 & n22916 ;
  assign n22918 = n22917 ^ n22915 ;
  assign n22920 = n22919 ^ n22918 ;
  assign n22921 = n22920 ^ n22205 ;
  assign n22922 = n22921 ^ n21429 ;
  assign n22909 = n22884 ^ n22874 ;
  assign n22910 = n22884 ^ n21071 ;
  assign n22911 = n22909 & n22910 ;
  assign n22912 = n22911 ^ n21071 ;
  assign n22913 = n22912 ^ n21112 ;
  assign n22923 = n22922 ^ n22913 ;
  assign n22925 = n22923 ^ x379 ;
  assign n22924 = n22923 ^ n22885 ;
  assign n22926 = n22925 ^ n22924 ;
  assign n22927 = n22890 & ~n22926 ;
  assign n22928 = n22927 ^ n22925 ;
  assign n22966 = n21885 ^ n21865 ;
  assign n22962 = n22241 ^ n22205 ;
  assign n22961 = n22919 ^ n22241 ;
  assign n22963 = n22962 ^ n22961 ;
  assign n22964 = n22918 & n22963 ;
  assign n22965 = n22964 ^ n22962 ;
  assign n22967 = n22966 ^ n22965 ;
  assign n22968 = n22967 ^ n22241 ;
  assign n22969 = n22968 ^ n21459 ;
  assign n22956 = n22922 ^ n22912 ;
  assign n22957 = n22922 ^ n21112 ;
  assign n22958 = n22956 & n22957 ;
  assign n22959 = n22958 ^ n21112 ;
  assign n22960 = n22959 ^ n21157 ;
  assign n22970 = n22969 ^ n22960 ;
  assign n22972 = n22970 ^ x378 ;
  assign n22971 = n22970 ^ n22923 ;
  assign n22973 = n22972 ^ n22971 ;
  assign n22974 = ~n22928 & n22973 ;
  assign n22975 = n22974 ^ n22972 ;
  assign n22929 = n22928 ^ x378 ;
  assign n22190 = n22151 & ~n22189 ;
  assign n22228 = n22227 ^ x367 ;
  assign n22229 = ~n22190 & n22228 ;
  assign n22267 = n22266 ^ x366 ;
  assign n22268 = ~n22229 & n22267 ;
  assign n22303 = n22302 ^ x365 ;
  assign n22304 = n22268 & n22303 ;
  assign n22320 = n22319 ^ x364 ;
  assign n22321 = n22304 & n22320 ;
  assign n22342 = n22341 ^ x363 ;
  assign n22343 = n22321 & ~n22342 ;
  assign n22363 = n22362 ^ x362 ;
  assign n22364 = ~n22343 & n22363 ;
  assign n22383 = n22382 ^ x361 ;
  assign n22384 = n22364 & ~n22383 ;
  assign n22405 = n22404 ^ x360 ;
  assign n22406 = ~n22384 & ~n22405 ;
  assign n22425 = n22424 ^ x375 ;
  assign n22426 = n22425 ^ n22421 ;
  assign n22434 = ~n22406 & n22426 ;
  assign n22456 = n22455 ^ x374 ;
  assign n22474 = ~n22434 & ~n22456 ;
  assign n22493 = n22492 ^ x373 ;
  assign n22510 = ~n22474 & ~n22493 ;
  assign n22527 = n22526 ^ x372 ;
  assign n22549 = n22510 & ~n22527 ;
  assign n22569 = n22568 ^ x371 ;
  assign n22590 = n22549 & ~n22569 ;
  assign n22610 = n22609 ^ x370 ;
  assign n22631 = ~n22590 & n22610 ;
  assign n22651 = n22650 ^ x369 ;
  assign n22672 = n22631 & n22651 ;
  assign n22692 = n22691 ^ x368 ;
  assign n22713 = ~n22672 & ~n22692 ;
  assign n22732 = n22731 ^ x383 ;
  assign n22733 = n22732 ^ n22728 ;
  assign n22753 = n22713 & n22733 ;
  assign n22774 = n22773 ^ x382 ;
  assign n22795 = ~n22753 & n22774 ;
  assign n22815 = n22814 ^ x381 ;
  assign n22836 = ~n22795 & n22815 ;
  assign n22856 = n22855 ^ x380 ;
  assign n22870 = n22836 & ~n22856 ;
  assign n22891 = n22890 ^ x379 ;
  assign n22930 = ~n22870 & ~n22891 ;
  assign n22977 = ~n22929 & ~n22930 ;
  assign n23012 = n22977 ^ n22970 ;
  assign n23013 = n22975 & ~n23012 ;
  assign n23010 = n22977 ^ n22975 ;
  assign n23011 = x377 & ~n23010 ;
  assign n23014 = n23013 ^ n23011 ;
  assign n23002 = n22966 ^ n22241 ;
  assign n23003 = n22965 & ~n23002 ;
  assign n22999 = n21906 ^ n21886 ;
  assign n23000 = n22999 ^ n22281 ;
  assign n23001 = n23000 ^ n22966 ;
  assign n23004 = n23003 ^ n23001 ;
  assign n23005 = n23004 ^ n22281 ;
  assign n23006 = n23005 ^ n21485 ;
  assign n23007 = n23006 ^ n21198 ;
  assign n22998 = n21157 ^ x376 ;
  assign n23008 = n23007 ^ n22998 ;
  assign n22995 = n22969 ^ n22959 ;
  assign n22996 = n22969 ^ n21157 ;
  assign n22997 = n22995 & n22996 ;
  assign n23009 = n23008 ^ n22997 ;
  assign n23015 = n23014 ^ n23009 ;
  assign n23058 = n23015 ^ n22391 ;
  assign n22892 = n22891 ^ n22870 ;
  assign n22932 = n22892 ^ n22334 ;
  assign n22432 = n21984 ^ n21951 ;
  assign n21930 = n21929 ^ n21928 ;
  assign n22427 = n22426 ^ n22406 ;
  assign n22431 = n21930 & n22427 ;
  assign n22433 = n22432 ^ n22431 ;
  assign n22468 = n21997 ^ n21983 ;
  assign n22457 = n22456 ^ n22434 ;
  assign n22469 = n22468 ^ n22457 ;
  assign n22470 = n22469 ^ n22431 ;
  assign n22471 = n22470 ^ n22468 ;
  assign n22472 = n22433 & n22471 ;
  assign n22473 = n22472 ^ n22469 ;
  assign n22503 = n21999 ^ n21515 ;
  assign n22504 = n22503 ^ n22019 ;
  assign n22494 = n22493 ^ n22474 ;
  assign n22506 = n22504 ^ n22494 ;
  assign n22505 = n22504 ^ n22468 ;
  assign n22507 = n22506 ^ n22505 ;
  assign n22508 = n22473 & ~n22507 ;
  assign n22509 = n22508 ^ n22505 ;
  assign n22542 = n22036 ^ n21512 ;
  assign n22543 = n22542 ^ n22061 ;
  assign n22545 = n22543 ^ n22504 ;
  assign n22528 = n22527 ^ n22510 ;
  assign n22544 = n22543 ^ n22528 ;
  assign n22546 = n22545 ^ n22544 ;
  assign n22547 = n22509 & n22546 ;
  assign n22548 = n22547 ^ n22545 ;
  assign n22584 = n22115 ^ n22097 ;
  assign n22570 = n22569 ^ n22549 ;
  assign n22586 = n22584 ^ n22570 ;
  assign n22585 = n22584 ^ n22543 ;
  assign n22587 = n22586 ^ n22585 ;
  assign n22588 = n22548 & n22587 ;
  assign n22589 = n22588 ^ n22585 ;
  assign n22624 = n22117 ^ n21580 ;
  assign n22625 = n22624 ^ n22137 ;
  assign n22627 = n22625 ^ n22584 ;
  assign n22611 = n22610 ^ n22590 ;
  assign n22626 = n22625 ^ n22611 ;
  assign n22628 = n22627 ^ n22626 ;
  assign n22629 = n22589 & ~n22628 ;
  assign n22630 = n22629 ^ n22627 ;
  assign n22665 = n22154 ^ n21594 ;
  assign n22666 = n22665 ^ n22176 ;
  assign n22652 = n22651 ^ n22631 ;
  assign n22668 = n22666 ^ n22652 ;
  assign n22667 = n22666 ^ n22625 ;
  assign n22669 = n22668 ^ n22667 ;
  assign n22670 = n22630 & n22669 ;
  assign n22671 = n22670 ^ n22667 ;
  assign n22706 = n22193 ^ n21633 ;
  assign n22707 = n22706 ^ n22215 ;
  assign n22693 = n22692 ^ n22672 ;
  assign n22709 = n22707 ^ n22693 ;
  assign n22708 = n22707 ^ n22666 ;
  assign n22710 = n22709 ^ n22708 ;
  assign n22711 = ~n22671 & n22710 ;
  assign n22712 = n22711 ^ n22708 ;
  assign n22747 = n22269 ^ n22251 ;
  assign n22734 = n22733 ^ n22713 ;
  assign n22749 = n22747 ^ n22734 ;
  assign n22748 = n22747 ^ n22707 ;
  assign n22750 = n22749 ^ n22748 ;
  assign n22751 = ~n22712 & ~n22750 ;
  assign n22752 = n22751 ^ n22748 ;
  assign n22788 = n22271 ^ n21677 ;
  assign n22789 = n22788 ^ n22290 ;
  assign n22791 = n22789 ^ n22747 ;
  assign n22775 = n22774 ^ n22753 ;
  assign n22790 = n22789 ^ n22775 ;
  assign n22792 = n22791 ^ n22790 ;
  assign n22793 = n22752 & ~n22792 ;
  assign n22794 = n22793 ^ n22791 ;
  assign n22829 = n21700 ^ n21608 ;
  assign n22830 = n22829 ^ n22311 ;
  assign n22832 = n22830 ^ n22789 ;
  assign n22816 = n22815 ^ n22795 ;
  assign n22831 = n22830 ^ n22816 ;
  assign n22833 = n22832 ^ n22831 ;
  assign n22834 = ~n22794 & ~n22833 ;
  assign n22835 = n22834 ^ n22832 ;
  assign n22857 = n22856 ^ n22836 ;
  assign n22893 = n22857 ^ n22830 ;
  assign n22894 = n22835 & ~n22893 ;
  assign n22895 = n22894 ^ n22830 ;
  assign n22933 = n22895 ^ n22892 ;
  assign n22934 = n22932 & n22933 ;
  assign n22935 = n22934 ^ n22334 ;
  assign n22931 = n22930 ^ n22929 ;
  assign n22949 = n22935 ^ n22931 ;
  assign n22950 = n22375 ^ n21767 ;
  assign n22951 = n22950 ^ n22354 ;
  assign n22952 = n22951 ^ n22931 ;
  assign n22953 = n22952 ^ n22950 ;
  assign n22954 = n22949 & n22953 ;
  assign n22955 = n22954 ^ n22951 ;
  assign n22976 = n22975 ^ x377 ;
  assign n22978 = n22977 ^ n22976 ;
  assign n23016 = n22978 ^ n22950 ;
  assign n23017 = ~n22955 & n23016 ;
  assign n23018 = n23017 ^ n22978 ;
  assign n23059 = n23018 ^ n23015 ;
  assign n23060 = n23058 & ~n23059 ;
  assign n23061 = n23060 ^ n22391 ;
  assign n23056 = n21955 ^ x359 ;
  assign n23115 = n23061 ^ n23056 ;
  assign n23116 = n23061 ^ n22413 ;
  assign n23117 = ~n23115 & ~n23116 ;
  assign n23118 = n23117 ^ n22413 ;
  assign n23201 = n23120 ^ n23118 ;
  assign n23202 = n21995 ^ n21961 ;
  assign n23203 = n23202 ^ n21961 ;
  assign n23204 = n23203 ^ n23202 ;
  assign n23205 = n23204 ^ n23118 ;
  assign n23206 = ~n23201 & ~n23205 ;
  assign n23207 = n23206 ^ n23203 ;
  assign n23208 = n22515 ^ n21873 ;
  assign n23210 = n23208 ^ n22482 ;
  assign n23209 = n23208 ^ n23202 ;
  assign n23211 = n23210 ^ n23209 ;
  assign n23212 = n23207 & ~n23211 ;
  assign n23213 = n23212 ^ n23210 ;
  assign n23214 = n22073 ^ n22033 ;
  assign n23217 = n23214 ^ n23208 ;
  assign n23215 = n22032 ^ n21996 ;
  assign n23216 = n23215 ^ n23214 ;
  assign n23218 = n23217 ^ n23216 ;
  assign n23219 = ~n23213 & n23218 ;
  assign n23220 = n23219 ^ n23217 ;
  assign n23222 = n22597 ^ n22556 ;
  assign n23221 = n23214 ^ n22597 ;
  assign n23223 = n23222 ^ n23221 ;
  assign n23224 = ~n23220 & n23223 ;
  assign n23225 = n23224 ^ n23222 ;
  assign n23228 = n22638 ^ n22597 ;
  assign n23226 = n22113 ^ n22074 ;
  assign n23227 = n23226 ^ n22638 ;
  assign n23229 = n23228 ^ n23227 ;
  assign n23230 = n23225 & ~n23229 ;
  assign n23231 = n23230 ^ n23228 ;
  assign n23234 = n22683 ^ n22638 ;
  assign n23232 = n22150 ^ n22114 ;
  assign n23233 = n23232 ^ n22683 ;
  assign n23235 = n23234 ^ n23233 ;
  assign n23236 = n23231 & n23235 ;
  assign n23237 = n23236 ^ n23234 ;
  assign n23290 = n23238 ^ n23237 ;
  assign n23291 = n23290 ^ n22684 ;
  assign n23284 = n23232 ^ n23231 ;
  assign n23285 = n23284 ^ n22639 ;
  assign n23278 = n23226 ^ n23225 ;
  assign n23279 = n23278 ^ n22598 ;
  assign n23272 = n23220 ^ n22556 ;
  assign n23273 = n23272 ^ n22557 ;
  assign n23266 = n23215 ^ n23213 ;
  assign n23267 = n23266 ^ n22515 ;
  assign n23256 = n23207 ^ n22482 ;
  assign n23257 = n23256 ^ n22483 ;
  assign n23258 = n23257 ^ n21844 ;
  assign n23019 = n23018 ^ n22391 ;
  assign n23020 = n23019 ^ n23015 ;
  assign n23021 = n23020 ^ n22392 ;
  assign n22529 = n22528 ^ n22509 ;
  assign n22530 = n22529 ^ n22020 ;
  assign n22573 = n22530 ^ n21445 ;
  assign n22495 = n22494 ^ n22473 ;
  assign n22496 = n22495 ^ n21987 ;
  assign n22458 = n22457 ^ n22433 ;
  assign n22459 = n22458 ^ n21953 ;
  assign n22429 = n22427 ^ n21411 ;
  assign n22430 = n21412 & n22429 ;
  assign n22460 = n22459 ^ n22430 ;
  assign n22464 = n22430 ^ n21414 ;
  assign n22465 = n22460 & ~n22464 ;
  assign n22466 = n22465 ^ n21414 ;
  assign n22531 = n22496 ^ n22466 ;
  assign n22532 = n22496 ^ n21416 ;
  assign n22533 = n22531 & n22532 ;
  assign n22534 = n22533 ^ n21416 ;
  assign n22574 = n22534 ^ n22530 ;
  assign n22575 = ~n22573 & n22574 ;
  assign n22576 = n22575 ^ n21445 ;
  assign n22577 = n22576 ^ n21474 ;
  assign n22571 = n22570 ^ n22548 ;
  assign n22572 = n22571 ^ n22062 ;
  assign n22614 = n22576 ^ n22572 ;
  assign n22615 = ~n22577 & n22614 ;
  assign n22616 = n22615 ^ n21474 ;
  assign n22617 = n22616 ^ n21504 ;
  assign n22612 = n22611 ^ n22589 ;
  assign n22613 = n22612 ^ n22101 ;
  assign n22655 = n22616 ^ n22613 ;
  assign n22656 = n22617 & ~n22655 ;
  assign n22657 = n22656 ^ n21504 ;
  assign n22658 = n22657 ^ n21573 ;
  assign n22653 = n22652 ^ n22630 ;
  assign n22654 = n22653 ^ n22138 ;
  assign n22696 = n22657 ^ n22654 ;
  assign n22697 = n22658 & n22696 ;
  assign n22698 = n22697 ^ n21573 ;
  assign n22699 = n22698 ^ n21588 ;
  assign n22694 = n22693 ^ n22671 ;
  assign n22695 = n22694 ^ n22177 ;
  assign n22737 = n22698 ^ n22695 ;
  assign n22738 = n22699 & ~n22737 ;
  assign n22739 = n22738 ^ n21588 ;
  assign n22740 = n22739 ^ n21627 ;
  assign n22735 = n22734 ^ n22712 ;
  assign n22736 = n22735 ^ n22216 ;
  assign n22778 = n22739 ^ n22736 ;
  assign n22779 = ~n22740 & n22778 ;
  assign n22780 = n22779 ^ n21627 ;
  assign n22781 = n22780 ^ n21652 ;
  assign n22776 = n22775 ^ n22752 ;
  assign n22777 = n22776 ^ n22255 ;
  assign n22819 = n22780 ^ n22777 ;
  assign n22820 = n22781 & n22819 ;
  assign n22821 = n22820 ^ n21652 ;
  assign n22822 = n22821 ^ n21670 ;
  assign n22817 = n22816 ^ n22794 ;
  assign n22818 = n22817 ^ n22291 ;
  assign n22860 = n22821 ^ n22818 ;
  assign n22861 = ~n22822 & n22860 ;
  assign n22862 = n22861 ^ n21670 ;
  assign n22863 = n22862 ^ n21693 ;
  assign n22858 = n22857 ^ n22835 ;
  assign n22859 = n22858 ^ n22312 ;
  assign n22899 = n22862 ^ n22859 ;
  assign n22900 = ~n22863 & ~n22899 ;
  assign n22901 = n22900 ^ n21693 ;
  assign n22902 = n22901 ^ n21715 ;
  assign n22896 = n22895 ^ n22334 ;
  assign n22897 = n22896 ^ n22892 ;
  assign n22898 = n22897 ^ n22335 ;
  assign n22939 = n22901 ^ n22898 ;
  assign n22940 = n22902 & ~n22939 ;
  assign n22941 = n22940 ^ n21715 ;
  assign n22942 = n22941 ^ n21738 ;
  assign n22936 = n22935 ^ n22354 ;
  assign n22937 = n22936 ^ n22931 ;
  assign n22938 = n22937 ^ n22355 ;
  assign n22981 = n22941 ^ n22938 ;
  assign n22982 = ~n22942 & ~n22981 ;
  assign n22983 = n22982 ^ n21738 ;
  assign n22984 = n22983 ^ n21760 ;
  assign n22979 = n22978 ^ n22955 ;
  assign n22980 = n22979 ^ n22375 ;
  assign n22991 = n22983 ^ n22980 ;
  assign n22992 = n22984 & ~n22991 ;
  assign n22993 = n22992 ^ n21760 ;
  assign n23055 = n23021 ^ n22993 ;
  assign n23057 = n23056 ^ n22413 ;
  assign n23062 = n23061 ^ n23057 ;
  assign n23063 = n23062 ^ n22414 ;
  assign n23064 = n23063 ^ n21781 ;
  assign n23065 = n23064 ^ n22993 ;
  assign n23066 = n23065 ^ n23063 ;
  assign n23067 = ~n23055 & n23066 ;
  assign n23068 = n23067 ^ n23064 ;
  assign n23119 = n23118 ^ n21961 ;
  assign n23121 = n23120 ^ n23119 ;
  assign n23122 = n23121 ^ n22443 ;
  assign n23124 = n23122 ^ n21808 ;
  assign n23123 = n23122 ^ n23063 ;
  assign n23125 = n23124 ^ n23123 ;
  assign n23126 = ~n23068 & n23125 ;
  assign n23127 = n23126 ^ n23124 ;
  assign n23260 = n23257 ^ n21822 ;
  assign n23259 = n23257 ^ n23122 ;
  assign n23261 = n23260 ^ n23259 ;
  assign n23262 = n23127 & ~n23261 ;
  assign n23263 = n23262 ^ n23260 ;
  assign n23264 = ~n23258 & n23263 ;
  assign n23265 = n23264 ^ n21844 ;
  assign n23268 = n23267 ^ n23265 ;
  assign n23269 = n23267 ^ n21866 ;
  assign n23270 = n23268 & n23269 ;
  assign n23271 = n23270 ^ n21866 ;
  assign n23274 = n23273 ^ n23271 ;
  assign n23275 = n23273 ^ n21887 ;
  assign n23276 = ~n23274 & ~n23275 ;
  assign n23277 = n23276 ^ n21887 ;
  assign n23280 = n23279 ^ n23277 ;
  assign n23281 = n23279 ^ n21911 ;
  assign n23282 = ~n23280 & n23281 ;
  assign n23283 = n23282 ^ n21911 ;
  assign n23286 = n23285 ^ n23283 ;
  assign n23287 = n23285 ^ n21273 ;
  assign n23288 = n23286 & ~n23287 ;
  assign n23289 = n23288 ^ n21273 ;
  assign n23292 = n23291 ^ n23289 ;
  assign n23240 = n22720 ^ n22683 ;
  assign n23239 = n23238 ^ n22720 ;
  assign n23241 = n23240 ^ n23239 ;
  assign n23242 = n23237 & ~n23241 ;
  assign n23243 = n23242 ^ n23240 ;
  assign n23199 = n22228 ^ n22190 ;
  assign n23293 = n23243 ^ n23199 ;
  assign n23294 = n23293 ^ n22721 ;
  assign n23295 = n23294 ^ n21294 ;
  assign n23296 = n23295 ^ n23294 ;
  assign n23297 = n23296 ^ n23289 ;
  assign n23298 = ~n23292 & ~n23297 ;
  assign n23299 = n23298 ^ n23295 ;
  assign n23415 = n23299 ^ n21316 ;
  assign n23371 = n23289 ^ n21294 ;
  assign n23372 = n23371 ^ n23291 ;
  assign n23373 = n23372 ^ x464 ;
  assign n22462 = x455 & ~n22429 ;
  assign n22461 = n22460 ^ n21414 ;
  assign n22463 = n22462 ^ n22461 ;
  assign n22467 = n22466 ^ n21416 ;
  assign n22497 = n22496 ^ n22467 ;
  assign n22498 = n22497 ^ x454 ;
  assign n22499 = n22498 ^ n22461 ;
  assign n22500 = n22499 ^ n22497 ;
  assign n22501 = ~n22463 & n22500 ;
  assign n22502 = n22501 ^ n22498 ;
  assign n22535 = n22534 ^ n21445 ;
  assign n22536 = n22535 ^ n22530 ;
  assign n22538 = n22536 ^ x453 ;
  assign n22537 = n22536 ^ n22497 ;
  assign n22539 = n22538 ^ n22537 ;
  assign n22540 = n22502 & ~n22539 ;
  assign n22541 = n22540 ^ n22538 ;
  assign n22578 = n22577 ^ n22572 ;
  assign n22580 = n22578 ^ x452 ;
  assign n22579 = n22578 ^ n22536 ;
  assign n22581 = n22580 ^ n22579 ;
  assign n22582 = n22541 & ~n22581 ;
  assign n22583 = n22582 ^ n22580 ;
  assign n22618 = n22617 ^ n22613 ;
  assign n22620 = n22618 ^ x451 ;
  assign n22619 = n22618 ^ n22578 ;
  assign n22621 = n22620 ^ n22619 ;
  assign n22622 = ~n22583 & n22621 ;
  assign n22623 = n22622 ^ n22620 ;
  assign n22659 = n22658 ^ n22654 ;
  assign n22661 = n22659 ^ x450 ;
  assign n22660 = n22659 ^ n22618 ;
  assign n22662 = n22661 ^ n22660 ;
  assign n22663 = n22623 & ~n22662 ;
  assign n22664 = n22663 ^ n22661 ;
  assign n22700 = n22699 ^ n22695 ;
  assign n22702 = n22700 ^ x449 ;
  assign n22701 = n22700 ^ n22659 ;
  assign n22703 = n22702 ^ n22701 ;
  assign n22704 = ~n22664 & n22703 ;
  assign n22705 = n22704 ^ n22702 ;
  assign n22741 = n22740 ^ n22736 ;
  assign n22743 = n22741 ^ x448 ;
  assign n22742 = n22741 ^ n22700 ;
  assign n22744 = n22743 ^ n22742 ;
  assign n22745 = n22705 & ~n22744 ;
  assign n22746 = n22745 ^ n22743 ;
  assign n22782 = n22781 ^ n22777 ;
  assign n22784 = n22782 ^ x463 ;
  assign n22783 = n22782 ^ n22741 ;
  assign n22785 = n22784 ^ n22783 ;
  assign n22786 = n22746 & ~n22785 ;
  assign n22787 = n22786 ^ n22784 ;
  assign n22823 = n22822 ^ n22818 ;
  assign n22825 = n22823 ^ x462 ;
  assign n22824 = n22823 ^ n22782 ;
  assign n22826 = n22825 ^ n22824 ;
  assign n22827 = n22787 & ~n22826 ;
  assign n22828 = n22827 ^ n22825 ;
  assign n22864 = n22863 ^ n22859 ;
  assign n22866 = n22864 ^ x461 ;
  assign n22865 = n22864 ^ n22823 ;
  assign n22867 = n22866 ^ n22865 ;
  assign n22868 = ~n22828 & n22867 ;
  assign n22869 = n22868 ^ n22866 ;
  assign n22903 = n22902 ^ n22898 ;
  assign n22905 = n22903 ^ x460 ;
  assign n22904 = n22903 ^ n22864 ;
  assign n22906 = n22905 ^ n22904 ;
  assign n22907 = ~n22869 & n22906 ;
  assign n22908 = n22907 ^ n22905 ;
  assign n22943 = n22942 ^ n22938 ;
  assign n22945 = n22943 ^ x459 ;
  assign n22944 = n22943 ^ n22903 ;
  assign n22946 = n22945 ^ n22944 ;
  assign n22947 = ~n22908 & n22946 ;
  assign n22948 = n22947 ^ n22945 ;
  assign n22985 = n22984 ^ n22980 ;
  assign n22987 = n22985 ^ x458 ;
  assign n22986 = n22985 ^ n22943 ;
  assign n22988 = n22987 ^ n22986 ;
  assign n22989 = n22948 & ~n22988 ;
  assign n22990 = n22989 ^ n22987 ;
  assign n22994 = n22993 ^ n21781 ;
  assign n23022 = n23021 ^ n22994 ;
  assign n23024 = n23022 ^ x457 ;
  assign n23023 = n23022 ^ n22985 ;
  assign n23025 = n23024 ^ n23023 ;
  assign n23026 = n22990 & ~n23025 ;
  assign n23027 = n23026 ^ n23024 ;
  assign n23070 = n23022 ^ x456 ;
  assign n23071 = n23027 & ~n23070 ;
  assign n23072 = n23071 ^ x456 ;
  assign n23069 = n23068 ^ n21808 ;
  assign n23114 = n23072 ^ n23069 ;
  assign n23128 = n23127 ^ n21822 ;
  assign n23129 = n23128 ^ x471 ;
  assign n23130 = n23129 ^ n23069 ;
  assign n23131 = n23130 ^ n23128 ;
  assign n23132 = n23114 & ~n23131 ;
  assign n23133 = n23132 ^ n23129 ;
  assign n23374 = n23263 ^ n21844 ;
  assign n23376 = n23374 ^ x470 ;
  assign n23375 = n23374 ^ n23128 ;
  assign n23377 = n23376 ^ n23375 ;
  assign n23378 = ~n23133 & n23377 ;
  assign n23379 = n23378 ^ n23376 ;
  assign n23380 = n23265 ^ n21866 ;
  assign n23381 = n23380 ^ n23267 ;
  assign n23383 = n23381 ^ x469 ;
  assign n23382 = n23381 ^ n23374 ;
  assign n23384 = n23383 ^ n23382 ;
  assign n23385 = ~n23379 & n23384 ;
  assign n23386 = n23385 ^ n23383 ;
  assign n23387 = n23271 ^ n21887 ;
  assign n23388 = n23387 ^ n23273 ;
  assign n23390 = n23388 ^ x468 ;
  assign n23389 = n23388 ^ n23381 ;
  assign n23391 = n23390 ^ n23389 ;
  assign n23392 = n23386 & ~n23391 ;
  assign n23393 = n23392 ^ n23390 ;
  assign n23394 = n23277 ^ n21911 ;
  assign n23395 = n23394 ^ n23279 ;
  assign n23397 = n23395 ^ x467 ;
  assign n23396 = n23395 ^ n23388 ;
  assign n23398 = n23397 ^ n23396 ;
  assign n23399 = n23393 & ~n23398 ;
  assign n23400 = n23399 ^ n23397 ;
  assign n23401 = n23283 ^ n21273 ;
  assign n23402 = n23401 ^ n23285 ;
  assign n23404 = n23402 ^ x466 ;
  assign n23403 = n23402 ^ n23395 ;
  assign n23405 = n23404 ^ n23403 ;
  assign n23406 = n23400 & ~n23405 ;
  assign n23407 = n23406 ^ n23404 ;
  assign n23409 = n23372 ^ x465 ;
  assign n23408 = n23402 ^ n23372 ;
  assign n23410 = n23409 ^ n23408 ;
  assign n23411 = ~n23407 & n23410 ;
  assign n23412 = n23411 ^ n23409 ;
  assign n23413 = n23373 & ~n23412 ;
  assign n23414 = n23413 ^ x464 ;
  assign n23416 = n23415 ^ n23414 ;
  assign n23247 = n22761 ^ n22047 ;
  assign n23200 = n23199 ^ n22720 ;
  assign n23244 = n23200 & n23243 ;
  assign n23245 = n23244 ^ n22720 ;
  assign n23198 = n22267 ^ n22229 ;
  assign n23246 = n23245 ^ n23198 ;
  assign n23300 = n23247 ^ n23246 ;
  assign n23301 = n23300 ^ n22761 ;
  assign n23303 = n23301 ^ n21316 ;
  assign n23302 = n23301 ^ n23294 ;
  assign n23304 = n23303 ^ n23302 ;
  assign n23305 = ~n23299 & ~n23304 ;
  assign n23306 = n23305 ^ n23303 ;
  assign n23417 = n23306 ^ n22040 ;
  assign n23418 = n23417 ^ x479 ;
  assign n23419 = n23418 ^ n23414 ;
  assign n23420 = n23419 ^ n23417 ;
  assign n23421 = n23416 & n23420 ;
  assign n23422 = n23421 ^ n23418 ;
  assign n23252 = n22303 ^ n22268 ;
  assign n23250 = n23247 ^ n22802 ;
  assign n23248 = n23247 ^ n23245 ;
  assign n23249 = n23246 & n23248 ;
  assign n23251 = n23250 ^ n23249 ;
  assign n23253 = n23252 ^ n23251 ;
  assign n23254 = n23253 ^ n22803 ;
  assign n23308 = n23254 ^ n22040 ;
  assign n23307 = n23301 ^ n23254 ;
  assign n23309 = n23308 ^ n23307 ;
  assign n23310 = ~n23306 & ~n23309 ;
  assign n23311 = n23310 ^ n23308 ;
  assign n23423 = n23311 ^ n22076 ;
  assign n23425 = n23423 ^ x478 ;
  assign n23424 = n23423 ^ n23417 ;
  assign n23426 = n23425 ^ n23424 ;
  assign n23427 = ~n23422 & n23426 ;
  assign n23428 = n23427 ^ n23425 ;
  assign n23255 = n23254 ^ n22076 ;
  assign n23312 = n23255 & n23311 ;
  assign n23313 = n23312 ^ n22076 ;
  assign n23429 = n23313 ^ n21379 ;
  assign n23319 = n22320 ^ n22304 ;
  assign n23315 = n22847 ^ n22802 ;
  assign n23314 = n23252 ^ n22847 ;
  assign n23316 = n23315 ^ n23314 ;
  assign n23317 = ~n23251 & ~n23316 ;
  assign n23318 = n23317 ^ n23315 ;
  assign n23320 = n23319 ^ n23318 ;
  assign n23321 = n23320 ^ n22848 ;
  assign n23430 = n23429 ^ n23321 ;
  assign n23432 = n23430 ^ x477 ;
  assign n23431 = n23430 ^ n23423 ;
  assign n23433 = n23432 ^ n23431 ;
  assign n23434 = ~n23428 & n23433 ;
  assign n23435 = n23434 ^ n23432 ;
  assign n23322 = n23321 ^ n23313 ;
  assign n23323 = n23321 ^ n21379 ;
  assign n23324 = ~n23322 & n23323 ;
  assign n23325 = n23324 ^ n21379 ;
  assign n23436 = n23325 ^ n21401 ;
  assign n23331 = n22342 ^ n22321 ;
  assign n23327 = n22882 ^ n22847 ;
  assign n23326 = n23319 ^ n22882 ;
  assign n23328 = n23327 ^ n23326 ;
  assign n23329 = ~n23318 & n23328 ;
  assign n23330 = n23329 ^ n23327 ;
  assign n23332 = n23331 ^ n23330 ;
  assign n23333 = n23332 ^ n22883 ;
  assign n23437 = n23436 ^ n23333 ;
  assign n23439 = n23437 ^ x476 ;
  assign n23438 = n23437 ^ n23430 ;
  assign n23440 = n23439 ^ n23438 ;
  assign n23441 = n23435 & ~n23440 ;
  assign n23442 = n23441 ^ n23439 ;
  assign n23334 = n23333 ^ n23325 ;
  assign n23335 = n23333 ^ n21401 ;
  assign n23336 = n23334 & ~n23335 ;
  assign n23337 = n23336 ^ n21401 ;
  assign n23443 = n23337 ^ n21429 ;
  assign n23343 = n22363 ^ n22343 ;
  assign n23339 = n22920 ^ n22882 ;
  assign n23338 = n23331 ^ n22920 ;
  assign n23340 = n23339 ^ n23338 ;
  assign n23341 = n23330 & ~n23340 ;
  assign n23342 = n23341 ^ n23339 ;
  assign n23344 = n23343 ^ n23342 ;
  assign n23345 = n23344 ^ n22921 ;
  assign n23444 = n23443 ^ n23345 ;
  assign n23446 = n23444 ^ x475 ;
  assign n23445 = n23444 ^ n23437 ;
  assign n23447 = n23446 ^ n23445 ;
  assign n23448 = ~n23442 & n23447 ;
  assign n23449 = n23448 ^ n23446 ;
  assign n23346 = n23345 ^ n23337 ;
  assign n23347 = n23345 ^ n21429 ;
  assign n23348 = ~n23346 & n23347 ;
  assign n23349 = n23348 ^ n21429 ;
  assign n23450 = n23349 ^ n21459 ;
  assign n23355 = n22383 ^ n22364 ;
  assign n23351 = n22967 ^ n22920 ;
  assign n23350 = n23343 ^ n22967 ;
  assign n23352 = n23351 ^ n23350 ;
  assign n23353 = ~n23342 & ~n23352 ;
  assign n23354 = n23353 ^ n23351 ;
  assign n23356 = n23355 ^ n23354 ;
  assign n23357 = n23356 ^ n22968 ;
  assign n23451 = n23450 ^ n23357 ;
  assign n23453 = n23451 ^ x474 ;
  assign n23452 = n23451 ^ n23444 ;
  assign n23454 = n23453 ^ n23452 ;
  assign n23455 = n23449 & ~n23454 ;
  assign n23456 = n23455 ^ n23453 ;
  assign n23490 = n23456 ^ x473 ;
  assign n23458 = n23422 ^ x478 ;
  assign n23459 = n23400 ^ x466 ;
  assign n23460 = n23393 ^ x467 ;
  assign n23461 = n23386 ^ x468 ;
  assign n23462 = n23379 ^ x469 ;
  assign n23028 = n23027 ^ x456 ;
  assign n23029 = n22990 ^ x457 ;
  assign n23030 = n22948 ^ x458 ;
  assign n23031 = n22908 ^ x459 ;
  assign n23032 = n22869 ^ x460 ;
  assign n23033 = n22828 ^ x461 ;
  assign n23034 = n22787 ^ x462 ;
  assign n23035 = n22502 ^ x453 ;
  assign n23036 = n22541 ^ x452 ;
  assign n23037 = n23035 & n23036 ;
  assign n23038 = n22583 ^ x451 ;
  assign n23039 = ~n23037 & n23038 ;
  assign n23040 = n22623 ^ x450 ;
  assign n23041 = n23039 & ~n23040 ;
  assign n23042 = n22664 ^ x449 ;
  assign n23043 = n23041 & n23042 ;
  assign n23044 = n22705 ^ x448 ;
  assign n23045 = n23043 & ~n23044 ;
  assign n23046 = n22746 ^ x463 ;
  assign n23047 = n23045 & ~n23046 ;
  assign n23048 = ~n23034 & n23047 ;
  assign n23049 = n23033 & n23048 ;
  assign n23050 = ~n23032 & ~n23049 ;
  assign n23051 = ~n23031 & n23050 ;
  assign n23052 = n23030 & n23051 ;
  assign n23053 = ~n23029 & ~n23052 ;
  assign n23054 = ~n23028 & n23053 ;
  assign n23073 = n23072 ^ x471 ;
  assign n23074 = n23073 ^ n23069 ;
  assign n23113 = ~n23054 & n23074 ;
  assign n23134 = n23133 ^ x470 ;
  assign n23463 = ~n23113 & n23134 ;
  assign n23464 = ~n23462 & ~n23463 ;
  assign n23465 = ~n23461 & ~n23464 ;
  assign n23466 = ~n23460 & n23465 ;
  assign n23467 = n23459 & ~n23466 ;
  assign n23468 = n23407 ^ x465 ;
  assign n23469 = n23467 & ~n23468 ;
  assign n23470 = n23412 ^ x464 ;
  assign n23471 = n23469 & ~n23470 ;
  assign n23472 = n23414 ^ x479 ;
  assign n23473 = n23472 ^ n23415 ;
  assign n23474 = n23471 & n23473 ;
  assign n23475 = n23458 & ~n23474 ;
  assign n23476 = n23428 ^ x477 ;
  assign n23477 = ~n23475 & ~n23476 ;
  assign n23478 = n23435 ^ x476 ;
  assign n23479 = n23477 & n23478 ;
  assign n23480 = n23442 ^ x475 ;
  assign n23481 = n23479 & ~n23480 ;
  assign n23482 = n23449 ^ x474 ;
  assign n23483 = n23481 & n23482 ;
  assign n23491 = n23490 ^ n23483 ;
  assign n23492 = n23491 ^ n23278 ;
  assign n23493 = n23482 ^ n23481 ;
  assign n23494 = n23493 ^ n23272 ;
  assign n23495 = n23480 ^ n23479 ;
  assign n23496 = n23495 ^ n23266 ;
  assign n23497 = n23478 ^ n23477 ;
  assign n23498 = n23497 ^ n23256 ;
  assign n23499 = n23476 ^ n23475 ;
  assign n23500 = n23499 ^ n23121 ;
  assign n23502 = n23470 ^ n23469 ;
  assign n23503 = n23502 ^ n22979 ;
  assign n23504 = n23468 ^ n23467 ;
  assign n23505 = n23504 ^ n22937 ;
  assign n23525 = n23466 ^ n23459 ;
  assign n23516 = n23464 ^ n23461 ;
  assign n23135 = n23134 ^ n23113 ;
  assign n23103 = n23053 ^ n23028 ;
  assign n23094 = n23051 ^ n23030 ;
  assign n23085 = n23049 ^ n23032 ;
  assign n23080 = n23048 ^ n23033 ;
  assign n22428 = n22427 ^ n21930 ;
  assign n23078 = n23047 ^ n23034 ;
  assign n23079 = n22428 & ~n23078 ;
  assign n23081 = n23080 ^ n23079 ;
  assign n23082 = n23080 ^ n22458 ;
  assign n23083 = ~n23081 & ~n23082 ;
  assign n23084 = n23083 ^ n22458 ;
  assign n23086 = n23085 ^ n23084 ;
  assign n23087 = n23085 ^ n22495 ;
  assign n23088 = ~n23086 & n23087 ;
  assign n23089 = n23088 ^ n22495 ;
  assign n23077 = n23050 ^ n23031 ;
  assign n23090 = n23089 ^ n23077 ;
  assign n23091 = n23089 ^ n22529 ;
  assign n23092 = n23090 & ~n23091 ;
  assign n23093 = n23092 ^ n22529 ;
  assign n23095 = n23094 ^ n23093 ;
  assign n23096 = n23094 ^ n22571 ;
  assign n23097 = n23095 & ~n23096 ;
  assign n23098 = n23097 ^ n22571 ;
  assign n23076 = n23052 ^ n23029 ;
  assign n23099 = n23098 ^ n23076 ;
  assign n23100 = n23098 ^ n22612 ;
  assign n23101 = ~n23099 & ~n23100 ;
  assign n23102 = n23101 ^ n22612 ;
  assign n23104 = n23103 ^ n23102 ;
  assign n23105 = n23103 ^ n22653 ;
  assign n23106 = ~n23104 & ~n23105 ;
  assign n23107 = n23106 ^ n22653 ;
  assign n23075 = n23074 ^ n23054 ;
  assign n23108 = n23107 ^ n23075 ;
  assign n23109 = n23107 ^ n22694 ;
  assign n23110 = ~n23108 & n23109 ;
  assign n23111 = n23110 ^ n22694 ;
  assign n23508 = n23135 ^ n23111 ;
  assign n23509 = n23135 ^ n22735 ;
  assign n23510 = n23508 & ~n23509 ;
  assign n23511 = n23510 ^ n22735 ;
  assign n23507 = n23463 ^ n23462 ;
  assign n23512 = n23511 ^ n23507 ;
  assign n23513 = n23511 ^ n22776 ;
  assign n23514 = n23512 & ~n23513 ;
  assign n23515 = n23514 ^ n22776 ;
  assign n23517 = n23516 ^ n23515 ;
  assign n23518 = n23516 ^ n22817 ;
  assign n23519 = n23517 & ~n23518 ;
  assign n23520 = n23519 ^ n22817 ;
  assign n23506 = n23465 ^ n23460 ;
  assign n23521 = n23520 ^ n23506 ;
  assign n23522 = n23520 ^ n22858 ;
  assign n23523 = ~n23521 & ~n23522 ;
  assign n23524 = n23523 ^ n22858 ;
  assign n23526 = n23525 ^ n23524 ;
  assign n23527 = n23525 ^ n22897 ;
  assign n23528 = ~n23526 & ~n23527 ;
  assign n23529 = n23528 ^ n22897 ;
  assign n23530 = n23529 ^ n23504 ;
  assign n23531 = n23505 & n23530 ;
  assign n23532 = n23531 ^ n22937 ;
  assign n23533 = n23532 ^ n23502 ;
  assign n23534 = ~n23503 & ~n23533 ;
  assign n23535 = n23534 ^ n22979 ;
  assign n23536 = n23535 ^ n23020 ;
  assign n23537 = n23473 ^ n23471 ;
  assign n23538 = n23537 ^ n23535 ;
  assign n23539 = n23536 & ~n23538 ;
  assign n23540 = n23539 ^ n23020 ;
  assign n23501 = n23474 ^ n23458 ;
  assign n23541 = n23540 ^ n23501 ;
  assign n23542 = n23499 ^ n23062 ;
  assign n23543 = n23542 ^ n23501 ;
  assign n23544 = n23543 ^ n23499 ;
  assign n23545 = ~n23541 & ~n23544 ;
  assign n23546 = n23545 ^ n23542 ;
  assign n23547 = n23500 & n23546 ;
  assign n23548 = n23547 ^ n23121 ;
  assign n23549 = n23548 ^ n23497 ;
  assign n23550 = ~n23498 & ~n23549 ;
  assign n23551 = n23550 ^ n23256 ;
  assign n23552 = n23551 ^ n23495 ;
  assign n23553 = ~n23496 & ~n23552 ;
  assign n23554 = n23553 ^ n23266 ;
  assign n23555 = n23554 ^ n23493 ;
  assign n23556 = ~n23494 & ~n23555 ;
  assign n23557 = n23556 ^ n23272 ;
  assign n23558 = n23557 ^ n23491 ;
  assign n23559 = ~n23492 & ~n23558 ;
  assign n23560 = n23559 ^ n23278 ;
  assign n23484 = n23483 ^ n23451 ;
  assign n23487 = ~n23456 & n23484 ;
  assign n23457 = n23456 ^ n23451 ;
  assign n23485 = n23484 ^ n23457 ;
  assign n23486 = x473 & n23485 ;
  assign n23488 = n23487 ^ n23486 ;
  assign n23365 = n23355 ^ n22967 ;
  assign n23366 = n23354 & n23365 ;
  assign n23363 = n22405 ^ n22384 ;
  assign n23362 = n23355 ^ n23004 ;
  assign n23364 = n23363 ^ n23362 ;
  assign n23367 = n23366 ^ n23364 ;
  assign n23368 = n23367 ^ n23006 ;
  assign n23361 = n21459 ^ x472 ;
  assign n23369 = n23368 ^ n23361 ;
  assign n23358 = n23357 ^ n23349 ;
  assign n23359 = n23357 ^ n21459 ;
  assign n23360 = ~n23358 & ~n23359 ;
  assign n23370 = n23369 ^ n23360 ;
  assign n23489 = n23488 ^ n23370 ;
  assign n23561 = n23560 ^ n23489 ;
  assign n23571 = n23561 ^ n22638 ;
  assign n23572 = n23571 ^ n21938 ;
  assign n23573 = n23558 ^ n22597 ;
  assign n23574 = n23573 ^ n21915 ;
  assign n23575 = n23555 ^ n22556 ;
  assign n23576 = n23575 ^ n21894 ;
  assign n23577 = n23552 ^ n23208 ;
  assign n23578 = n23577 ^ n21873 ;
  assign n23579 = n23549 ^ n22482 ;
  assign n23580 = n23579 ^ n21851 ;
  assign n23582 = n23546 ^ n22443 ;
  assign n23642 = n23541 ^ n22413 ;
  assign n23583 = n23538 ^ n22391 ;
  assign n23584 = n23583 ^ n21788 ;
  assign n23585 = n23533 ^ n22950 ;
  assign n23586 = n23585 ^ n21767 ;
  assign n23587 = n23530 ^ n22354 ;
  assign n23588 = n23587 ^ n21745 ;
  assign n23589 = n23526 ^ n22334 ;
  assign n23590 = n23589 ^ n21722 ;
  assign n23625 = n23521 ^ n22830 ;
  assign n23620 = n23517 ^ n22789 ;
  assign n23615 = n23512 ^ n22747 ;
  assign n23610 = n23508 ^ n22707 ;
  assign n23605 = n23108 ^ n22666 ;
  assign n23600 = n23104 ^ n22625 ;
  assign n23595 = n23099 ^ n22584 ;
  assign n23172 = n23095 ^ n22543 ;
  assign n23160 = n23090 ^ n22504 ;
  assign n23148 = n23086 ^ n22468 ;
  assign n23139 = n23081 ^ n22432 ;
  assign n23137 = n23078 ^ n21928 ;
  assign n23138 = ~n21929 & ~n23137 ;
  assign n23140 = n23139 ^ n23138 ;
  assign n23144 = n23138 ^ n21520 ;
  assign n23145 = n23140 & ~n23144 ;
  assign n23146 = n23145 ^ n21520 ;
  assign n23155 = n23148 ^ n23146 ;
  assign n23156 = n23148 ^ n21526 ;
  assign n23157 = n23155 & ~n23156 ;
  assign n23158 = n23157 ^ n21526 ;
  assign n23167 = n23160 ^ n23158 ;
  assign n23168 = n23160 ^ n21515 ;
  assign n23169 = ~n23167 & n23168 ;
  assign n23170 = n23169 ^ n21515 ;
  assign n23591 = n23172 ^ n23170 ;
  assign n23592 = n23172 ^ n21512 ;
  assign n23593 = ~n23591 & n23592 ;
  assign n23594 = n23593 ^ n21512 ;
  assign n23596 = n23595 ^ n23594 ;
  assign n23597 = n23595 ^ n21510 ;
  assign n23598 = n23596 & n23597 ;
  assign n23599 = n23598 ^ n21510 ;
  assign n23601 = n23600 ^ n23599 ;
  assign n23602 = n23600 ^ n21580 ;
  assign n23603 = ~n23601 & n23602 ;
  assign n23604 = n23603 ^ n21580 ;
  assign n23606 = n23605 ^ n23604 ;
  assign n23607 = n23605 ^ n21594 ;
  assign n23608 = n23606 & ~n23607 ;
  assign n23609 = n23608 ^ n21594 ;
  assign n23611 = n23610 ^ n23609 ;
  assign n23612 = n23610 ^ n21633 ;
  assign n23613 = n23611 & ~n23612 ;
  assign n23614 = n23613 ^ n21633 ;
  assign n23616 = n23615 ^ n23614 ;
  assign n23617 = n23615 ^ n21655 ;
  assign n23618 = n23616 & ~n23617 ;
  assign n23619 = n23618 ^ n21655 ;
  assign n23621 = n23620 ^ n23619 ;
  assign n23622 = n23620 ^ n21677 ;
  assign n23623 = ~n23621 & ~n23622 ;
  assign n23624 = n23623 ^ n21677 ;
  assign n23626 = n23625 ^ n23624 ;
  assign n23627 = n23625 ^ n21700 ;
  assign n23628 = ~n23626 & ~n23627 ;
  assign n23629 = n23628 ^ n21700 ;
  assign n23630 = n23629 ^ n23589 ;
  assign n23631 = ~n23590 & ~n23630 ;
  assign n23632 = n23631 ^ n21722 ;
  assign n23633 = n23632 ^ n23587 ;
  assign n23634 = ~n23588 & n23633 ;
  assign n23635 = n23634 ^ n21745 ;
  assign n23636 = n23635 ^ n23585 ;
  assign n23637 = n23586 & ~n23636 ;
  assign n23638 = n23637 ^ n21767 ;
  assign n23639 = n23638 ^ n23583 ;
  assign n23640 = n23584 & ~n23639 ;
  assign n23641 = n23640 ^ n21788 ;
  assign n23643 = n23642 ^ n23641 ;
  assign n23644 = n23120 ^ n21815 ;
  assign n23645 = n23644 ^ n23546 ;
  assign n23646 = n23645 ^ n23120 ;
  assign n23647 = n23646 ^ n23641 ;
  assign n23648 = n23647 ^ n23546 ;
  assign n23649 = n23643 & n23648 ;
  assign n23650 = n23649 ^ n23645 ;
  assign n23651 = n23582 & ~n23650 ;
  assign n23581 = n23579 ^ n21829 ;
  assign n23652 = n23651 ^ n23581 ;
  assign n23653 = n23580 & ~n23652 ;
  assign n23654 = n23653 ^ n21851 ;
  assign n23655 = n23654 ^ n23577 ;
  assign n23656 = ~n23578 & n23655 ;
  assign n23657 = n23656 ^ n21873 ;
  assign n23658 = n23657 ^ n23575 ;
  assign n23659 = n23576 & n23658 ;
  assign n23660 = n23659 ^ n21894 ;
  assign n23661 = n23660 ^ n23573 ;
  assign n23662 = n23574 & ~n23661 ;
  assign n23663 = n23662 ^ n21915 ;
  assign n23664 = n23663 ^ n23571 ;
  assign n23665 = n23572 & ~n23664 ;
  assign n23666 = n23665 ^ n21938 ;
  assign n23684 = n23666 ^ n21971 ;
  assign n23567 = n22429 ^ x455 ;
  assign n23562 = n23290 ^ n23284 ;
  assign n23563 = n23562 ^ n23290 ;
  assign n23564 = n23563 ^ n23489 ;
  assign n23565 = ~n23561 & ~n23564 ;
  assign n23566 = n23565 ^ n23562 ;
  assign n23568 = n23567 ^ n23566 ;
  assign n23569 = n23568 ^ n23290 ;
  assign n23570 = n23569 ^ n22683 ;
  assign n23685 = n23684 ^ n23570 ;
  assign n23686 = n23685 ^ x48 ;
  assign n23767 = n23641 ^ n21815 ;
  assign n23768 = n23767 ^ n23642 ;
  assign n23687 = n23638 ^ n21788 ;
  assign n23688 = n23687 ^ n23583 ;
  assign n23689 = n23688 ^ x40 ;
  assign n23142 = x39 & n23137 ;
  assign n23141 = n23140 ^ n21520 ;
  assign n23143 = n23142 ^ n23141 ;
  assign n23147 = n23146 ^ n21526 ;
  assign n23149 = n23148 ^ n23147 ;
  assign n23150 = n23149 ^ x38 ;
  assign n23151 = n23150 ^ n23141 ;
  assign n23152 = n23151 ^ n23149 ;
  assign n23153 = ~n23143 & n23152 ;
  assign n23154 = n23153 ^ n23150 ;
  assign n23159 = n23158 ^ n21515 ;
  assign n23161 = n23160 ^ n23159 ;
  assign n23163 = n23161 ^ x37 ;
  assign n23162 = n23161 ^ n23149 ;
  assign n23164 = n23163 ^ n23162 ;
  assign n23165 = ~n23154 & n23164 ;
  assign n23166 = n23165 ^ n23163 ;
  assign n23171 = n23170 ^ n21512 ;
  assign n23173 = n23172 ^ n23171 ;
  assign n23175 = n23173 ^ x36 ;
  assign n23174 = n23173 ^ n23161 ;
  assign n23176 = n23175 ^ n23174 ;
  assign n23177 = n23166 & ~n23176 ;
  assign n23178 = n23177 ^ n23175 ;
  assign n23690 = n23594 ^ n21510 ;
  assign n23691 = n23690 ^ n23595 ;
  assign n23693 = n23691 ^ x35 ;
  assign n23692 = n23691 ^ n23173 ;
  assign n23694 = n23693 ^ n23692 ;
  assign n23695 = n23178 & ~n23694 ;
  assign n23696 = n23695 ^ n23693 ;
  assign n23697 = n23599 ^ n21580 ;
  assign n23698 = n23697 ^ n23600 ;
  assign n23700 = n23698 ^ x34 ;
  assign n23699 = n23698 ^ n23691 ;
  assign n23701 = n23700 ^ n23699 ;
  assign n23702 = n23696 & ~n23701 ;
  assign n23703 = n23702 ^ n23700 ;
  assign n23704 = n23604 ^ n21594 ;
  assign n23705 = n23704 ^ n23605 ;
  assign n23707 = n23705 ^ x33 ;
  assign n23706 = n23705 ^ n23698 ;
  assign n23708 = n23707 ^ n23706 ;
  assign n23709 = ~n23703 & n23708 ;
  assign n23710 = n23709 ^ n23707 ;
  assign n23711 = n23609 ^ n21633 ;
  assign n23712 = n23711 ^ n23610 ;
  assign n23714 = n23712 ^ x32 ;
  assign n23713 = n23712 ^ n23705 ;
  assign n23715 = n23714 ^ n23713 ;
  assign n23716 = n23710 & ~n23715 ;
  assign n23717 = n23716 ^ n23714 ;
  assign n23718 = n23614 ^ n21655 ;
  assign n23719 = n23718 ^ n23615 ;
  assign n23721 = n23719 ^ x47 ;
  assign n23720 = n23719 ^ n23712 ;
  assign n23722 = n23721 ^ n23720 ;
  assign n23723 = n23717 & ~n23722 ;
  assign n23724 = n23723 ^ n23721 ;
  assign n23725 = n23619 ^ n21677 ;
  assign n23726 = n23725 ^ n23620 ;
  assign n23728 = n23726 ^ x46 ;
  assign n23727 = n23726 ^ n23719 ;
  assign n23729 = n23728 ^ n23727 ;
  assign n23730 = n23724 & ~n23729 ;
  assign n23731 = n23730 ^ n23728 ;
  assign n23732 = n23624 ^ n21700 ;
  assign n23733 = n23732 ^ n23625 ;
  assign n23735 = n23733 ^ x45 ;
  assign n23734 = n23733 ^ n23726 ;
  assign n23736 = n23735 ^ n23734 ;
  assign n23737 = n23731 & ~n23736 ;
  assign n23738 = n23737 ^ n23735 ;
  assign n23739 = n23629 ^ n21722 ;
  assign n23740 = n23739 ^ n23589 ;
  assign n23742 = n23740 ^ x44 ;
  assign n23741 = n23740 ^ n23733 ;
  assign n23743 = n23742 ^ n23741 ;
  assign n23744 = ~n23738 & n23743 ;
  assign n23745 = n23744 ^ n23742 ;
  assign n23746 = n23632 ^ n21745 ;
  assign n23747 = n23746 ^ n23587 ;
  assign n23749 = n23747 ^ x43 ;
  assign n23748 = n23747 ^ n23740 ;
  assign n23750 = n23749 ^ n23748 ;
  assign n23751 = n23745 & ~n23750 ;
  assign n23752 = n23751 ^ n23749 ;
  assign n23753 = n23635 ^ n21767 ;
  assign n23754 = n23753 ^ n23585 ;
  assign n23756 = n23754 ^ x42 ;
  assign n23755 = n23754 ^ n23747 ;
  assign n23757 = n23756 ^ n23755 ;
  assign n23758 = ~n23752 & n23757 ;
  assign n23759 = n23758 ^ n23756 ;
  assign n23761 = n23688 ^ x41 ;
  assign n23760 = n23754 ^ n23688 ;
  assign n23762 = n23761 ^ n23760 ;
  assign n23763 = n23759 & ~n23762 ;
  assign n23764 = n23763 ^ n23761 ;
  assign n23765 = ~n23689 & n23764 ;
  assign n23766 = n23765 ^ x40 ;
  assign n23769 = n23768 ^ n23766 ;
  assign n23770 = n23650 ^ n21829 ;
  assign n23771 = n23770 ^ x55 ;
  assign n23772 = n23771 ^ n23766 ;
  assign n23773 = n23772 ^ n23770 ;
  assign n23774 = ~n23769 & n23773 ;
  assign n23775 = n23774 ^ n23771 ;
  assign n23776 = n23652 ^ n21851 ;
  assign n23778 = n23776 ^ x54 ;
  assign n23777 = n23776 ^ n23770 ;
  assign n23779 = n23778 ^ n23777 ;
  assign n23780 = n23775 & ~n23779 ;
  assign n23781 = n23780 ^ n23778 ;
  assign n23782 = n23654 ^ n21873 ;
  assign n23783 = n23782 ^ n23577 ;
  assign n23785 = n23783 ^ x53 ;
  assign n23784 = n23783 ^ n23776 ;
  assign n23786 = n23785 ^ n23784 ;
  assign n23787 = n23781 & ~n23786 ;
  assign n23788 = n23787 ^ n23785 ;
  assign n23789 = n23657 ^ n21894 ;
  assign n23790 = n23789 ^ n23575 ;
  assign n23792 = n23790 ^ x52 ;
  assign n23791 = n23790 ^ n23783 ;
  assign n23793 = n23792 ^ n23791 ;
  assign n23794 = ~n23788 & n23793 ;
  assign n23795 = n23794 ^ n23792 ;
  assign n23796 = n23660 ^ n21915 ;
  assign n23797 = n23796 ^ n23573 ;
  assign n23799 = n23797 ^ x51 ;
  assign n23798 = n23797 ^ n23790 ;
  assign n23800 = n23799 ^ n23798 ;
  assign n23801 = n23795 & ~n23800 ;
  assign n23802 = n23801 ^ n23799 ;
  assign n23803 = n23663 ^ n21938 ;
  assign n23804 = n23803 ^ n23571 ;
  assign n23806 = n23804 ^ x50 ;
  assign n23805 = n23804 ^ n23797 ;
  assign n23807 = n23806 ^ n23805 ;
  assign n23808 = ~n23802 & n23807 ;
  assign n23809 = n23808 ^ n23806 ;
  assign n23811 = n23685 ^ x49 ;
  assign n23810 = n23804 ^ n23685 ;
  assign n23812 = n23811 ^ n23810 ;
  assign n23813 = ~n23809 & n23812 ;
  assign n23814 = n23813 ^ n23811 ;
  assign n23815 = ~n23686 & n23814 ;
  assign n23816 = n23815 ^ x48 ;
  assign n23667 = n23666 ^ n23570 ;
  assign n23673 = n22462 ^ x454 ;
  assign n23674 = n23673 ^ n22461 ;
  assign n23669 = n23293 ^ n23290 ;
  assign n23668 = n23567 ^ n23293 ;
  assign n23670 = n23669 ^ n23668 ;
  assign n23671 = ~n23566 & n23670 ;
  assign n23672 = n23671 ^ n23669 ;
  assign n23675 = n23674 ^ n23672 ;
  assign n23676 = n23675 ^ n23293 ;
  assign n23677 = n23676 ^ n22720 ;
  assign n23678 = n23677 ^ n21971 ;
  assign n23679 = n23678 ^ n23570 ;
  assign n23680 = n23679 ^ n23677 ;
  assign n23681 = n23667 & ~n23680 ;
  assign n23682 = n23681 ^ n23678 ;
  assign n23683 = n23682 ^ n22015 ;
  assign n23817 = n23816 ^ n23683 ;
  assign n23824 = n23247 ^ n22015 ;
  assign n23819 = n23674 ^ n23293 ;
  assign n23820 = ~n23672 & n23819 ;
  assign n23821 = n23820 ^ n23293 ;
  assign n23822 = n23821 ^ n23035 ;
  assign n23825 = n23824 ^ n23822 ;
  assign n23818 = n23677 ^ n23247 ;
  assign n23823 = n23822 ^ n23818 ;
  assign n23826 = n23825 ^ n23823 ;
  assign n23827 = n23682 & ~n23826 ;
  assign n23828 = n23827 ^ n23825 ;
  assign n23829 = n23828 ^ n22047 ;
  assign n23830 = n23829 ^ x63 ;
  assign n23831 = n23830 ^ n23683 ;
  assign n23832 = n23831 ^ n23829 ;
  assign n23833 = n23817 & ~n23832 ;
  assign n23834 = n23833 ^ n23830 ;
  assign n23846 = n23822 ^ n22761 ;
  assign n23847 = ~n23828 & n23846 ;
  assign n23841 = n23036 ^ n23035 ;
  assign n23835 = n23821 ^ n23300 ;
  assign n23836 = n23253 ^ n23035 ;
  assign n23837 = n23836 ^ n23253 ;
  assign n23838 = n23837 ^ n23821 ;
  assign n23839 = n23835 & n23838 ;
  assign n23840 = n23839 ^ n23836 ;
  assign n23842 = n23841 ^ n23840 ;
  assign n23843 = n23842 ^ n23253 ;
  assign n23844 = n23843 ^ n22802 ;
  assign n23845 = n23844 ^ n22047 ;
  assign n23848 = n23847 ^ n23845 ;
  assign n23849 = n23848 ^ n22083 ;
  assign n23851 = n23849 ^ x62 ;
  assign n23850 = n23849 ^ n23829 ;
  assign n23852 = n23851 ^ n23850 ;
  assign n23853 = ~n23834 & n23852 ;
  assign n23854 = n23853 ^ n23851 ;
  assign n23864 = n23038 ^ n23037 ;
  assign n23860 = n23320 ^ n23253 ;
  assign n23859 = n23841 ^ n23320 ;
  assign n23861 = n23860 ^ n23859 ;
  assign n23862 = ~n23840 & n23861 ;
  assign n23863 = n23862 ^ n23860 ;
  assign n23865 = n23864 ^ n23863 ;
  assign n23866 = n23865 ^ n23320 ;
  assign n23867 = n23866 ^ n22847 ;
  assign n23855 = n23844 ^ n22083 ;
  assign n23856 = ~n23848 & ~n23855 ;
  assign n23857 = n23856 ^ n22083 ;
  assign n23858 = n23857 ^ n22128 ;
  assign n23868 = n23867 ^ n23858 ;
  assign n23870 = n23868 ^ x61 ;
  assign n23869 = n23868 ^ n23849 ;
  assign n23871 = n23870 ^ n23869 ;
  assign n23872 = n23854 & ~n23871 ;
  assign n23873 = n23872 ^ n23870 ;
  assign n23879 = n23040 ^ n23039 ;
  assign n23881 = n23879 ^ n23320 ;
  assign n23880 = n23879 ^ n23864 ;
  assign n23882 = n23881 ^ n23880 ;
  assign n23883 = n23863 & n23882 ;
  assign n23884 = n23883 ^ n23881 ;
  assign n23885 = n23884 ^ n22882 ;
  assign n23874 = n23867 ^ n23857 ;
  assign n23875 = n23867 ^ n22128 ;
  assign n23876 = n23874 & n23875 ;
  assign n23877 = n23876 ^ n22128 ;
  assign n23878 = n23877 ^ n22166 ;
  assign n23886 = n23885 ^ n23878 ;
  assign n23888 = n23886 ^ x60 ;
  assign n23887 = n23886 ^ n23868 ;
  assign n23889 = n23888 ^ n23887 ;
  assign n23890 = n23873 & ~n23889 ;
  assign n23891 = n23890 ^ n23888 ;
  assign n23980 = n23891 ^ x59 ;
  assign n23931 = n23745 ^ x43 ;
  assign n23932 = n23738 ^ x44 ;
  assign n23179 = n23178 ^ x35 ;
  assign n23180 = n23154 ^ x37 ;
  assign n23181 = n23166 ^ x36 ;
  assign n23182 = n23180 & ~n23181 ;
  assign n23933 = ~n23179 & n23182 ;
  assign n23934 = n23696 ^ x34 ;
  assign n23935 = n23933 & ~n23934 ;
  assign n23936 = n23703 ^ x33 ;
  assign n23937 = ~n23935 & ~n23936 ;
  assign n23938 = n23710 ^ x32 ;
  assign n23939 = ~n23937 & ~n23938 ;
  assign n23940 = n23717 ^ x47 ;
  assign n23941 = n23939 & ~n23940 ;
  assign n23942 = n23724 ^ x46 ;
  assign n23943 = ~n23941 & n23942 ;
  assign n23944 = n23731 ^ x45 ;
  assign n23945 = ~n23943 & ~n23944 ;
  assign n23946 = ~n23932 & ~n23945 ;
  assign n23947 = ~n23931 & ~n23946 ;
  assign n23948 = n23752 ^ x42 ;
  assign n23949 = ~n23947 & ~n23948 ;
  assign n23950 = n23759 ^ x41 ;
  assign n23951 = n23949 & n23950 ;
  assign n23952 = n23764 ^ x40 ;
  assign n23953 = n23951 & n23952 ;
  assign n23954 = n23766 ^ x55 ;
  assign n23955 = n23954 ^ n23768 ;
  assign n23956 = ~n23953 & n23955 ;
  assign n23957 = n23775 ^ x54 ;
  assign n23958 = ~n23956 & n23957 ;
  assign n23959 = n23781 ^ x53 ;
  assign n23960 = n23958 & n23959 ;
  assign n23961 = n23788 ^ x52 ;
  assign n23962 = n23960 & ~n23961 ;
  assign n23963 = n23795 ^ x51 ;
  assign n23964 = n23962 & n23963 ;
  assign n23965 = n23802 ^ x50 ;
  assign n23966 = n23964 & ~n23965 ;
  assign n23967 = n23809 ^ x49 ;
  assign n23968 = ~n23966 & n23967 ;
  assign n23969 = n23814 ^ x48 ;
  assign n23970 = ~n23968 & n23969 ;
  assign n23971 = n23816 ^ x63 ;
  assign n23972 = n23971 ^ n23683 ;
  assign n23973 = ~n23970 & ~n23972 ;
  assign n23974 = n23834 ^ x62 ;
  assign n23975 = n23973 & n23974 ;
  assign n23976 = n23854 ^ x61 ;
  assign n23977 = ~n23975 & n23976 ;
  assign n23978 = n23873 ^ x60 ;
  assign n23979 = ~n23977 & ~n23978 ;
  assign n23987 = n23980 ^ n23979 ;
  assign n24192 = n23987 ^ n22427 ;
  assign n24193 = x135 & ~n24192 ;
  assign n24097 = n23987 ^ n22428 ;
  assign n24098 = n21930 & ~n24097 ;
  assign n24190 = n24098 ^ n22432 ;
  assign n23902 = n23042 ^ n23041 ;
  assign n23898 = n23344 ^ n23332 ;
  assign n23897 = n23879 ^ n23344 ;
  assign n23899 = n23898 ^ n23897 ;
  assign n23900 = ~n23884 & n23899 ;
  assign n23901 = n23900 ^ n23898 ;
  assign n23903 = n23902 ^ n23901 ;
  assign n23904 = n23903 ^ n23344 ;
  assign n23905 = n23904 ^ n22920 ;
  assign n23892 = n23885 ^ n23877 ;
  assign n23893 = n23885 ^ n22166 ;
  assign n23894 = ~n23892 & ~n23893 ;
  assign n23895 = n23894 ^ n22166 ;
  assign n23896 = n23895 ^ n22205 ;
  assign n23906 = n23905 ^ n23896 ;
  assign n23908 = n23906 ^ x59 ;
  assign n23907 = n23906 ^ n23886 ;
  assign n23909 = n23908 ^ n23907 ;
  assign n23910 = n23891 & ~n23909 ;
  assign n23911 = n23910 ^ n23908 ;
  assign n23982 = n23911 ^ x58 ;
  assign n23981 = n23979 & ~n23980 ;
  assign n23992 = n23982 ^ n23981 ;
  assign n23989 = n23079 ^ n22458 ;
  assign n23990 = n23989 ^ n23080 ;
  assign n23986 = n23078 ^ n22428 ;
  assign n23988 = ~n23986 & ~n23987 ;
  assign n23991 = n23990 ^ n23988 ;
  assign n24095 = n23992 ^ n23991 ;
  assign n24096 = n24095 ^ n23081 ;
  assign n24191 = n24190 ^ n24096 ;
  assign n24194 = n24193 ^ n24191 ;
  assign n24099 = n24098 ^ n24096 ;
  assign n23993 = n23992 ^ n23988 ;
  assign n23994 = ~n23991 & n23993 ;
  assign n23995 = n23994 ^ n23990 ;
  assign n23196 = n23084 ^ n22495 ;
  assign n23197 = n23196 ^ n23085 ;
  assign n23996 = n23995 ^ n23197 ;
  assign n23983 = ~n23981 & ~n23982 ;
  assign n23917 = n23044 ^ n23043 ;
  assign n23919 = n23917 ^ n23344 ;
  assign n23918 = n23917 ^ n23902 ;
  assign n23920 = n23919 ^ n23918 ;
  assign n23921 = n23901 & ~n23920 ;
  assign n23922 = n23921 ^ n23919 ;
  assign n23923 = n23922 ^ n22967 ;
  assign n23912 = n23905 ^ n23895 ;
  assign n23913 = n23905 ^ n22205 ;
  assign n23914 = n23912 & ~n23913 ;
  assign n23915 = n23914 ^ n22205 ;
  assign n23916 = n23915 ^ n22241 ;
  assign n23924 = n23923 ^ n23916 ;
  assign n23926 = n23924 ^ x58 ;
  assign n23925 = n23924 ^ n23906 ;
  assign n23927 = n23926 ^ n23925 ;
  assign n23928 = ~n23911 & n23927 ;
  assign n23929 = n23928 ^ n23926 ;
  assign n23930 = n23929 ^ x57 ;
  assign n23984 = n23983 ^ n23930 ;
  assign n24092 = n23996 ^ n23984 ;
  assign n24093 = n24092 ^ n23086 ;
  assign n24100 = n24093 ^ n22432 ;
  assign n24101 = n24100 ^ n24093 ;
  assign n24102 = n24101 ^ n24096 ;
  assign n24103 = ~n24099 & ~n24102 ;
  assign n24104 = n24103 ^ n24100 ;
  assign n24195 = n24104 ^ n22468 ;
  assign n24196 = n24195 ^ x134 ;
  assign n24197 = n24196 ^ n24191 ;
  assign n24198 = n24197 ^ n24195 ;
  assign n24199 = n24194 & ~n24198 ;
  assign n24200 = n24199 ^ n24196 ;
  assign n24017 = n23983 ^ n23924 ;
  assign n24020 = n23929 & ~n24017 ;
  assign n24016 = n23929 ^ n23924 ;
  assign n24018 = n24017 ^ n24016 ;
  assign n24019 = ~x57 & n24018 ;
  assign n24021 = n24020 ^ n24019 ;
  assign n24008 = n23917 ^ n23356 ;
  assign n24009 = n23922 & n24008 ;
  assign n24005 = n23367 ^ n23045 ;
  assign n24006 = n24005 ^ n23046 ;
  assign n24007 = n24006 ^ n23917 ;
  assign n24010 = n24009 ^ n24007 ;
  assign n24011 = n24010 ^ n23367 ;
  assign n24012 = n24011 ^ n23004 ;
  assign n24013 = n24012 ^ n22281 ;
  assign n24004 = n22241 ^ x56 ;
  assign n24014 = n24013 ^ n24004 ;
  assign n24001 = n23923 ^ n23915 ;
  assign n24002 = n23923 ^ n22241 ;
  assign n24003 = n24001 & n24002 ;
  assign n24015 = n24014 ^ n24003 ;
  assign n24022 = n24021 ^ n24015 ;
  assign n23998 = n23091 ^ n23077 ;
  assign n23999 = n23998 ^ n23984 ;
  assign n23985 = n23984 ^ n23197 ;
  assign n23997 = ~n23985 & ~n23996 ;
  assign n24000 = n23999 ^ n23997 ;
  assign n24108 = n24022 ^ n24000 ;
  assign n24109 = n24108 ^ n23090 ;
  assign n24094 = n24093 ^ n22468 ;
  assign n24105 = n24094 & n24104 ;
  assign n24106 = n24105 ^ n22468 ;
  assign n24107 = n24106 ^ n22504 ;
  assign n24201 = n24109 ^ n24107 ;
  assign n24203 = n24201 ^ x133 ;
  assign n24202 = n24201 ^ n24195 ;
  assign n24204 = n24203 ^ n24202 ;
  assign n24205 = n24200 & ~n24204 ;
  assign n24206 = n24205 ^ n24203 ;
  assign n24027 = n23137 ^ x39 ;
  assign n23193 = n23093 ^ n22571 ;
  assign n23194 = n23193 ^ n23094 ;
  assign n24025 = n24022 ^ n23194 ;
  assign n24023 = n24022 ^ n23998 ;
  assign n24024 = n24000 & ~n24023 ;
  assign n24026 = n24025 ^ n24024 ;
  assign n24114 = n24027 ^ n24026 ;
  assign n24115 = n24114 ^ n23095 ;
  assign n24110 = n24109 ^ n24106 ;
  assign n24111 = n24107 & ~n24110 ;
  assign n24112 = n24111 ^ n22504 ;
  assign n24113 = n24112 ^ n22543 ;
  assign n24207 = n24115 ^ n24113 ;
  assign n24209 = n24207 ^ x132 ;
  assign n24208 = n24207 ^ n24201 ;
  assign n24210 = n24209 ^ n24208 ;
  assign n24211 = ~n24206 & n24210 ;
  assign n24212 = n24211 ^ n24209 ;
  assign n24028 = n24027 ^ n23194 ;
  assign n24029 = ~n24026 & ~n24028 ;
  assign n23189 = n23100 ^ n23076 ;
  assign n23195 = n23194 ^ n23189 ;
  assign n24030 = n24029 ^ n23195 ;
  assign n23190 = n23142 ^ x38 ;
  assign n23191 = n23190 ^ n23141 ;
  assign n24120 = n24030 ^ n23191 ;
  assign n24121 = n24120 ^ n23099 ;
  assign n24116 = n24115 ^ n24112 ;
  assign n24117 = n24113 & ~n24116 ;
  assign n24118 = n24117 ^ n22543 ;
  assign n24119 = n24118 ^ n22584 ;
  assign n24213 = n24121 ^ n24119 ;
  assign n24215 = n24213 ^ x131 ;
  assign n24214 = n24213 ^ n24207 ;
  assign n24216 = n24215 ^ n24214 ;
  assign n24217 = ~n24212 & n24216 ;
  assign n24218 = n24217 ^ n24215 ;
  assign n24396 = n24218 ^ x130 ;
  assign n24397 = n24192 ^ x135 ;
  assign n24398 = n24193 ^ x134 ;
  assign n24399 = n24398 ^ n24191 ;
  assign n24400 = ~n24397 & ~n24399 ;
  assign n24401 = n24200 ^ x133 ;
  assign n24402 = n24400 & ~n24401 ;
  assign n24403 = n24206 ^ x132 ;
  assign n24404 = ~n24402 & ~n24403 ;
  assign n24405 = n24212 ^ x131 ;
  assign n24406 = ~n24404 & n24405 ;
  assign n24407 = ~n24396 & ~n24406 ;
  assign n24122 = n24121 ^ n24118 ;
  assign n24123 = n24119 & ~n24122 ;
  assign n24124 = n24123 ^ n22584 ;
  assign n24187 = n24124 ^ n22625 ;
  assign n24033 = n23102 ^ n22653 ;
  assign n24034 = n24033 ^ n23103 ;
  assign n24125 = n24034 ^ n23180 ;
  assign n23192 = n23191 ^ n23189 ;
  assign n24031 = ~n23192 & ~n24030 ;
  assign n24032 = n24031 ^ n23191 ;
  assign n24126 = n24125 ^ n24032 ;
  assign n24127 = n24126 ^ n23104 ;
  assign n24188 = n24187 ^ n24127 ;
  assign n24220 = n24188 ^ x130 ;
  assign n24219 = n24213 ^ n24188 ;
  assign n24221 = n24220 ^ n24219 ;
  assign n24222 = ~n24218 & n24221 ;
  assign n24223 = n24222 ^ n24220 ;
  assign n24408 = n24223 ^ x129 ;
  assign n24409 = ~n24407 & ~n24408 ;
  assign n24189 = n24188 ^ x129 ;
  assign n24224 = ~n24189 & n24223 ;
  assign n24225 = n24224 ^ x129 ;
  assign n24128 = n24127 ^ n24124 ;
  assign n24129 = n24127 ^ n22625 ;
  assign n24130 = n24128 & ~n24129 ;
  assign n24131 = n24130 ^ n22625 ;
  assign n24185 = n24131 ^ n22666 ;
  assign n24035 = n24034 ^ n24032 ;
  assign n23185 = n23109 ^ n23075 ;
  assign n24036 = n23185 ^ n23180 ;
  assign n24037 = n24036 ^ n23185 ;
  assign n24038 = n24037 ^ n24032 ;
  assign n24039 = ~n24035 & ~n24038 ;
  assign n24040 = n24039 ^ n24036 ;
  assign n23187 = n23181 ^ n23180 ;
  assign n24089 = n24040 ^ n23187 ;
  assign n24090 = n24089 ^ n23108 ;
  assign n24186 = n24185 ^ n24090 ;
  assign n24226 = n24225 ^ n24186 ;
  assign n24410 = n24226 ^ x128 ;
  assign n24411 = ~n24409 & n24410 ;
  assign n23188 = n23187 ^ n23185 ;
  assign n24041 = ~n23188 & ~n24040 ;
  assign n23112 = n23111 ^ n22735 ;
  assign n23136 = n23135 ^ n23112 ;
  assign n23186 = n23185 ^ n23136 ;
  assign n24042 = n24041 ^ n23186 ;
  assign n23183 = n23182 ^ n23179 ;
  assign n24136 = n24042 ^ n23183 ;
  assign n24137 = n24136 ^ n23508 ;
  assign n24091 = n24090 ^ n22666 ;
  assign n24132 = n24131 ^ n24090 ;
  assign n24133 = ~n24091 & ~n24132 ;
  assign n24134 = n24133 ^ n22666 ;
  assign n24135 = n24134 ^ n22707 ;
  assign n24227 = n24137 ^ n24135 ;
  assign n24228 = n24227 ^ x128 ;
  assign n24229 = n24228 ^ n24225 ;
  assign n24230 = n24229 ^ n24227 ;
  assign n24231 = n24226 & n24230 ;
  assign n24232 = n24231 ^ n24228 ;
  assign n24412 = n24232 ^ x143 ;
  assign n24413 = n24411 & ~n24412 ;
  assign n24047 = n23513 ^ n23507 ;
  assign n24045 = n23934 ^ n23933 ;
  assign n23184 = n23183 ^ n23136 ;
  assign n24043 = n23184 & n24042 ;
  assign n24044 = n24043 ^ n23183 ;
  assign n24046 = n24045 ^ n24044 ;
  assign n24142 = n24047 ^ n24046 ;
  assign n24143 = n24142 ^ n23512 ;
  assign n24138 = n24137 ^ n24134 ;
  assign n24139 = ~n24135 & ~n24138 ;
  assign n24140 = n24139 ^ n22707 ;
  assign n24141 = n24140 ^ n22747 ;
  assign n24233 = n24143 ^ n24141 ;
  assign n24235 = n24233 ^ x143 ;
  assign n24234 = n24233 ^ n24227 ;
  assign n24236 = n24235 ^ n24234 ;
  assign n24237 = ~n24232 & n24236 ;
  assign n24238 = n24237 ^ n24235 ;
  assign n24414 = n24238 ^ x142 ;
  assign n24415 = n24413 & n24414 ;
  assign n24057 = n23936 ^ n23935 ;
  assign n24050 = n23515 ^ n22817 ;
  assign n24051 = n24050 ^ n23516 ;
  assign n24052 = n24051 ^ n24047 ;
  assign n24048 = n24047 ^ n24044 ;
  assign n24049 = ~n24046 & ~n24048 ;
  assign n24053 = n24052 ^ n24049 ;
  assign n24148 = n24057 ^ n24053 ;
  assign n24149 = n24148 ^ n23517 ;
  assign n24144 = n24143 ^ n24140 ;
  assign n24145 = n24141 & n24144 ;
  assign n24146 = n24145 ^ n22747 ;
  assign n24147 = n24146 ^ n22789 ;
  assign n24239 = n24149 ^ n24147 ;
  assign n24241 = n24239 ^ x142 ;
  assign n24240 = n24239 ^ n24233 ;
  assign n24242 = n24241 ^ n24240 ;
  assign n24243 = n24238 & ~n24242 ;
  assign n24244 = n24243 ^ n24241 ;
  assign n24416 = n24244 ^ x141 ;
  assign n24417 = n24415 & n24416 ;
  assign n24061 = n23938 ^ n23937 ;
  assign n24054 = n23522 ^ n23506 ;
  assign n24055 = n24054 ^ n24051 ;
  assign n24056 = n24055 ^ n24054 ;
  assign n24058 = n24057 ^ n24056 ;
  assign n24059 = n24053 & ~n24058 ;
  assign n24060 = n24059 ^ n24055 ;
  assign n24154 = n24061 ^ n24060 ;
  assign n24155 = n24154 ^ n23521 ;
  assign n24150 = n24149 ^ n24146 ;
  assign n24151 = ~n24147 & ~n24150 ;
  assign n24152 = n24151 ^ n22789 ;
  assign n24153 = n24152 ^ n22830 ;
  assign n24245 = n24155 ^ n24153 ;
  assign n24247 = n24245 ^ x141 ;
  assign n24246 = n24245 ^ n24239 ;
  assign n24248 = n24247 ^ n24246 ;
  assign n24249 = n24244 & ~n24248 ;
  assign n24250 = n24249 ^ n24247 ;
  assign n24418 = n24250 ^ x140 ;
  assign n24419 = n24417 & ~n24418 ;
  assign n24069 = n23940 ^ n23939 ;
  assign n24062 = n23524 ^ n22897 ;
  assign n24063 = n24062 ^ n23525 ;
  assign n24065 = n24063 ^ n24054 ;
  assign n24064 = n24063 ^ n24061 ;
  assign n24066 = n24065 ^ n24064 ;
  assign n24067 = n24060 & n24066 ;
  assign n24068 = n24067 ^ n24065 ;
  assign n24160 = n24069 ^ n24068 ;
  assign n24161 = n24160 ^ n23526 ;
  assign n24156 = n24155 ^ n24152 ;
  assign n24157 = n24153 & n24156 ;
  assign n24158 = n24157 ^ n22830 ;
  assign n24159 = n24158 ^ n22334 ;
  assign n24251 = n24161 ^ n24159 ;
  assign n24253 = n24251 ^ x140 ;
  assign n24252 = n24251 ^ n24245 ;
  assign n24254 = n24253 ^ n24252 ;
  assign n24255 = ~n24250 & n24254 ;
  assign n24256 = n24255 ^ n24253 ;
  assign n24420 = n24256 ^ x139 ;
  assign n24421 = ~n24419 & ~n24420 ;
  assign n24077 = n23942 ^ n23941 ;
  assign n24070 = n23529 ^ n22937 ;
  assign n24071 = n24070 ^ n23504 ;
  assign n24073 = n24071 ^ n24063 ;
  assign n24072 = n24071 ^ n24069 ;
  assign n24074 = n24073 ^ n24072 ;
  assign n24075 = ~n24068 & n24074 ;
  assign n24076 = n24075 ^ n24073 ;
  assign n24166 = n24077 ^ n24076 ;
  assign n24167 = n24166 ^ n23530 ;
  assign n24162 = n24161 ^ n24158 ;
  assign n24163 = ~n24159 & n24162 ;
  assign n24164 = n24163 ^ n22334 ;
  assign n24165 = n24164 ^ n22354 ;
  assign n24257 = n24167 ^ n24165 ;
  assign n24259 = n24257 ^ x139 ;
  assign n24258 = n24257 ^ n24251 ;
  assign n24260 = n24259 ^ n24258 ;
  assign n24261 = n24256 & ~n24260 ;
  assign n24262 = n24261 ^ n24259 ;
  assign n24422 = n24262 ^ x138 ;
  assign n24423 = n24421 & n24422 ;
  assign n24168 = n24167 ^ n24164 ;
  assign n24169 = ~n24165 & n24168 ;
  assign n24170 = n24169 ^ n22354 ;
  assign n24263 = n24170 ^ n22950 ;
  assign n24085 = n23944 ^ n23943 ;
  assign n24078 = n23532 ^ n22979 ;
  assign n24079 = n24078 ^ n23502 ;
  assign n24081 = n24079 ^ n24071 ;
  assign n24080 = n24079 ^ n24077 ;
  assign n24082 = n24081 ^ n24080 ;
  assign n24083 = n24076 & ~n24082 ;
  assign n24084 = n24083 ^ n24081 ;
  assign n24086 = n24085 ^ n24084 ;
  assign n24087 = n24086 ^ n23533 ;
  assign n24264 = n24263 ^ n24087 ;
  assign n24266 = n24264 ^ x138 ;
  assign n24265 = n24264 ^ n24257 ;
  assign n24267 = n24266 ^ n24265 ;
  assign n24268 = ~n24262 & n24267 ;
  assign n24269 = n24268 ^ n24266 ;
  assign n24424 = n24269 ^ x137 ;
  assign n24425 = ~n24423 & ~n24424 ;
  assign n24180 = n23945 ^ n23932 ;
  assign n24177 = n24085 ^ n24079 ;
  assign n24178 = n24084 & ~n24177 ;
  assign n24175 = n23537 ^ n23536 ;
  assign n24176 = n24175 ^ n24079 ;
  assign n24179 = n24178 ^ n24176 ;
  assign n24181 = n24180 ^ n24179 ;
  assign n24182 = n24181 ^ n23538 ;
  assign n24088 = n24087 ^ n22950 ;
  assign n24171 = n24170 ^ n24087 ;
  assign n24172 = ~n24088 & n24171 ;
  assign n24173 = n24172 ^ n22950 ;
  assign n24174 = n24173 ^ n22391 ;
  assign n24183 = n24182 ^ n24174 ;
  assign n24271 = n24183 ^ x137 ;
  assign n24270 = n24264 ^ n24183 ;
  assign n24272 = n24271 ^ n24270 ;
  assign n24273 = ~n24269 & n24272 ;
  assign n24274 = n24273 ^ n24271 ;
  assign n24426 = n24274 ^ x136 ;
  assign n24427 = n24425 & n24426 ;
  assign n24184 = n24183 ^ x136 ;
  assign n24275 = ~n24184 & n24274 ;
  assign n24276 = n24275 ^ x136 ;
  assign n24428 = n24276 ^ x151 ;
  assign n24277 = n24182 ^ n24173 ;
  assign n24283 = n23946 ^ n23931 ;
  assign n24281 = n23501 ^ n23062 ;
  assign n24282 = n24281 ^ n23540 ;
  assign n24284 = n24283 ^ n24282 ;
  assign n24278 = n24180 ^ n24175 ;
  assign n24279 = ~n24179 & n24278 ;
  assign n24280 = n24279 ^ n24180 ;
  assign n24285 = n24284 ^ n24280 ;
  assign n24286 = n24285 ^ n23541 ;
  assign n24287 = n24286 ^ n22391 ;
  assign n24288 = n24287 ^ n24173 ;
  assign n24289 = n24288 ^ n24286 ;
  assign n24290 = ~n24277 & n24289 ;
  assign n24291 = n24290 ^ n24287 ;
  assign n24292 = n24291 ^ n22413 ;
  assign n24429 = n24428 ^ n24292 ;
  assign n24430 = ~n24427 & n24429 ;
  assign n24293 = n24292 ^ n24276 ;
  assign n24298 = n23948 ^ n23947 ;
  assign n24295 = n24282 ^ n24280 ;
  assign n24296 = n24284 & n24295 ;
  assign n24297 = n24296 ^ n24283 ;
  assign n24299 = n24298 ^ n24297 ;
  assign n24294 = n23546 ^ n23121 ;
  assign n24300 = n24299 ^ n24294 ;
  assign n24301 = n24300 ^ n23546 ;
  assign n24303 = n24301 ^ n22413 ;
  assign n24302 = n24301 ^ n24286 ;
  assign n24304 = n24303 ^ n24302 ;
  assign n24305 = ~n24291 & ~n24304 ;
  assign n24306 = n24305 ^ n24303 ;
  assign n24307 = n24306 ^ n23120 ;
  assign n24308 = n24307 ^ x151 ;
  assign n24309 = n24308 ^ n24276 ;
  assign n24310 = n24309 ^ n24307 ;
  assign n24311 = ~n24293 & n24310 ;
  assign n24312 = n24311 ^ n24308 ;
  assign n24431 = n24312 ^ x150 ;
  assign n24432 = ~n24430 & ~n24431 ;
  assign n24316 = n23548 ^ n23256 ;
  assign n24317 = n24316 ^ n23497 ;
  assign n24318 = n24317 ^ n24294 ;
  assign n24314 = n24297 ^ n24294 ;
  assign n24315 = n24299 & n24314 ;
  assign n24319 = n24318 ^ n24315 ;
  assign n24313 = n23950 ^ n23949 ;
  assign n24320 = n24319 ^ n24313 ;
  assign n24321 = n24320 ^ n23549 ;
  assign n24323 = n24321 ^ n23120 ;
  assign n24322 = n24321 ^ n24301 ;
  assign n24324 = n24323 ^ n24322 ;
  assign n24325 = ~n24306 & n24324 ;
  assign n24326 = n24325 ^ n24323 ;
  assign n24327 = n24326 ^ n22482 ;
  assign n24329 = n24327 ^ x150 ;
  assign n24328 = n24327 ^ n24307 ;
  assign n24330 = n24329 ^ n24328 ;
  assign n24331 = ~n24312 & n24330 ;
  assign n24332 = n24331 ^ n24329 ;
  assign n24433 = n24332 ^ x149 ;
  assign n24434 = n24432 & ~n24433 ;
  assign n24344 = n23952 ^ n23951 ;
  assign n24337 = n23551 ^ n23266 ;
  assign n24338 = n24337 ^ n23495 ;
  assign n24339 = n24338 ^ n24317 ;
  assign n24340 = n24339 ^ n24338 ;
  assign n24341 = n24340 ^ n24313 ;
  assign n24342 = n24319 & ~n24341 ;
  assign n24343 = n24342 ^ n24339 ;
  assign n24345 = n24344 ^ n24343 ;
  assign n24346 = n24345 ^ n23552 ;
  assign n24333 = n24321 ^ n22482 ;
  assign n24334 = n24326 & n24333 ;
  assign n24335 = n24334 ^ n22482 ;
  assign n24336 = n24335 ^ n23208 ;
  assign n24347 = n24346 ^ n24336 ;
  assign n24349 = n24347 ^ x149 ;
  assign n24348 = n24347 ^ n24327 ;
  assign n24350 = n24349 ^ n24348 ;
  assign n24351 = ~n24332 & n24350 ;
  assign n24352 = n24351 ^ n24349 ;
  assign n24435 = n24352 ^ x148 ;
  assign n24436 = n24434 & n24435 ;
  assign n24365 = n23955 ^ n23953 ;
  assign n24358 = n23554 ^ n23272 ;
  assign n24359 = n24358 ^ n23493 ;
  assign n24361 = n24359 ^ n24338 ;
  assign n24360 = n24359 ^ n24344 ;
  assign n24362 = n24361 ^ n24360 ;
  assign n24363 = ~n24343 & n24362 ;
  assign n24364 = n24363 ^ n24361 ;
  assign n24366 = n24365 ^ n24364 ;
  assign n24367 = n24366 ^ n23555 ;
  assign n24353 = n24346 ^ n23208 ;
  assign n24354 = n24346 ^ n24335 ;
  assign n24355 = n24353 & n24354 ;
  assign n24356 = n24355 ^ n23208 ;
  assign n24357 = n24356 ^ n22556 ;
  assign n24368 = n24367 ^ n24357 ;
  assign n24370 = n24368 ^ x148 ;
  assign n24369 = n24368 ^ n24347 ;
  assign n24371 = n24370 ^ n24369 ;
  assign n24372 = n24352 & ~n24371 ;
  assign n24373 = n24372 ^ n24370 ;
  assign n24437 = n24373 ^ x147 ;
  assign n24438 = n24436 & ~n24437 ;
  assign n24386 = n23957 ^ n23956 ;
  assign n24379 = n23557 ^ n23278 ;
  assign n24380 = n24379 ^ n23491 ;
  assign n24382 = n24380 ^ n24359 ;
  assign n24381 = n24380 ^ n24365 ;
  assign n24383 = n24382 ^ n24381 ;
  assign n24384 = ~n24364 & ~n24383 ;
  assign n24385 = n24384 ^ n24382 ;
  assign n24387 = n24386 ^ n24385 ;
  assign n24388 = n24387 ^ n23558 ;
  assign n24374 = n24367 ^ n22556 ;
  assign n24375 = n24367 ^ n24356 ;
  assign n24376 = n24374 & ~n24375 ;
  assign n24377 = n24376 ^ n22556 ;
  assign n24378 = n24377 ^ n22597 ;
  assign n24389 = n24388 ^ n24378 ;
  assign n24391 = n24389 ^ x147 ;
  assign n24390 = n24389 ^ n24368 ;
  assign n24392 = n24391 ^ n24390 ;
  assign n24393 = ~n24373 & n24392 ;
  assign n24394 = n24393 ^ n24391 ;
  assign n24395 = n24394 ^ x146 ;
  assign n24439 = n24438 ^ n24395 ;
  assign n24440 = n24439 ^ n23078 ;
  assign n24472 = x231 & ~n24440 ;
  assign n24467 = n24097 ^ n23078 ;
  assign n24468 = n24439 & n24467 ;
  assign n24465 = ~n24395 & ~n24438 ;
  assign n24455 = n23959 ^ n23958 ;
  assign n24448 = n23560 ^ n23284 ;
  assign n24449 = n24448 ^ n23489 ;
  assign n24451 = n24449 ^ n24380 ;
  assign n24450 = n24449 ^ n24386 ;
  assign n24452 = n24451 ^ n24450 ;
  assign n24453 = ~n24385 & ~n24452 ;
  assign n24454 = n24453 ^ n24451 ;
  assign n24456 = n24455 ^ n24454 ;
  assign n24457 = n24456 ^ n23561 ;
  assign n24443 = n24388 ^ n22597 ;
  assign n24444 = n24388 ^ n24377 ;
  assign n24445 = ~n24443 & n24444 ;
  assign n24446 = n24445 ^ n22597 ;
  assign n24447 = n24446 ^ n22638 ;
  assign n24458 = n24457 ^ n24447 ;
  assign n24460 = n24458 ^ x146 ;
  assign n24459 = n24458 ^ n24389 ;
  assign n24461 = n24460 ^ n24459 ;
  assign n24462 = n24394 & ~n24461 ;
  assign n24463 = n24462 ^ n24460 ;
  assign n24464 = n24463 ^ x145 ;
  assign n24466 = n24465 ^ n24464 ;
  assign n24469 = n24468 ^ n24466 ;
  assign n24470 = n24469 ^ n23990 ;
  assign n24441 = n22428 & n24440 ;
  assign n24442 = n24441 ^ n22458 ;
  assign n24471 = n24470 ^ n24442 ;
  assign n24473 = n24472 ^ n24471 ;
  assign n24499 = n24468 ^ n24095 ;
  assign n24500 = n24469 & n24499 ;
  assign n24501 = n24500 ^ n24095 ;
  assign n24497 = ~n24464 & ~n24465 ;
  assign n24485 = n24455 ^ n24449 ;
  assign n24486 = ~n24454 & ~n24485 ;
  assign n24484 = n24449 ^ n23568 ;
  assign n24487 = n24486 ^ n24484 ;
  assign n24483 = n23961 ^ n23960 ;
  assign n24488 = n24487 ^ n24483 ;
  assign n24489 = n24488 ^ n23569 ;
  assign n24478 = n24457 ^ n22638 ;
  assign n24479 = n24457 ^ n24446 ;
  assign n24480 = n24478 & ~n24479 ;
  assign n24481 = n24480 ^ n22638 ;
  assign n24482 = n24481 ^ n22683 ;
  assign n24490 = n24489 ^ n24482 ;
  assign n24492 = n24490 ^ x145 ;
  assign n24491 = n24490 ^ n24458 ;
  assign n24493 = n24492 ^ n24491 ;
  assign n24494 = ~n24463 & n24493 ;
  assign n24495 = n24494 ^ n24492 ;
  assign n24496 = n24495 ^ x144 ;
  assign n24498 = n24497 ^ n24496 ;
  assign n24502 = n24501 ^ n24498 ;
  assign n24503 = n24502 ^ n23197 ;
  assign n24474 = n24470 ^ n24441 ;
  assign n24475 = ~n24442 & ~n24474 ;
  assign n24476 = n24475 ^ n22458 ;
  assign n24477 = n24476 ^ n22495 ;
  assign n24504 = n24503 ^ n24477 ;
  assign n24505 = n24504 ^ x230 ;
  assign n24506 = n24505 ^ n24472 ;
  assign n24507 = n24506 ^ n24504 ;
  assign n24508 = n24473 & n24507 ;
  assign n24509 = n24508 ^ n24505 ;
  assign n24536 = n24496 & n24497 ;
  assign n24521 = n24489 ^ n24481 ;
  assign n24524 = n24483 ^ n23568 ;
  assign n24525 = n24487 & n24524 ;
  assign n24526 = n24525 ^ n23568 ;
  assign n24522 = n23963 ^ n23962 ;
  assign n24523 = n24522 ^ n23675 ;
  assign n24527 = n24526 ^ n24523 ;
  assign n24528 = n24527 ^ n23676 ;
  assign n24529 = n24528 ^ n22683 ;
  assign n24530 = n24529 ^ n24481 ;
  assign n24531 = n24530 ^ n24528 ;
  assign n24532 = n24521 & n24531 ;
  assign n24533 = n24532 ^ n24529 ;
  assign n24534 = n24533 ^ n22720 ;
  assign n24517 = n24490 ^ x144 ;
  assign n24518 = n24495 & ~n24517 ;
  assign n24519 = n24518 ^ x144 ;
  assign n24520 = n24519 ^ x159 ;
  assign n24535 = n24534 ^ n24520 ;
  assign n24537 = n24536 ^ n24535 ;
  assign n24514 = n24501 ^ n24092 ;
  assign n24515 = n24502 & n24514 ;
  assign n24516 = n24515 ^ n24092 ;
  assign n24538 = n24537 ^ n24516 ;
  assign n24539 = n24538 ^ n23998 ;
  assign n24510 = n24503 ^ n24476 ;
  assign n24511 = n24477 & n24510 ;
  assign n24512 = n24511 ^ n22495 ;
  assign n24513 = n24512 ^ n22529 ;
  assign n24540 = n24539 ^ n24513 ;
  assign n24542 = n24540 ^ x229 ;
  assign n24541 = n24540 ^ n24504 ;
  assign n24543 = n24542 ^ n24541 ;
  assign n24544 = ~n24509 & n24543 ;
  assign n24545 = n24544 ^ n24542 ;
  assign n24576 = n24535 & n24536 ;
  assign n24553 = n24534 ^ n24519 ;
  assign n24561 = n23965 ^ n23964 ;
  assign n24554 = n24526 ^ n24522 ;
  assign n24555 = n23822 ^ n23300 ;
  assign n24556 = n24555 ^ n23675 ;
  assign n24557 = n24556 ^ n24522 ;
  assign n24558 = n24557 ^ n24555 ;
  assign n24559 = n24554 & n24558 ;
  assign n24560 = n24559 ^ n24556 ;
  assign n24562 = n24561 ^ n24560 ;
  assign n24563 = n24562 ^ n23822 ;
  assign n24565 = n24563 ^ n22720 ;
  assign n24564 = n24563 ^ n24528 ;
  assign n24566 = n24565 ^ n24564 ;
  assign n24567 = n24533 & ~n24566 ;
  assign n24568 = n24567 ^ n24565 ;
  assign n24569 = n24568 ^ n23247 ;
  assign n24570 = n24569 ^ x159 ;
  assign n24571 = n24570 ^ n24519 ;
  assign n24572 = n24571 ^ n24569 ;
  assign n24573 = n24553 & n24572 ;
  assign n24574 = n24573 ^ n24570 ;
  assign n24575 = n24574 ^ x158 ;
  assign n24577 = n24576 ^ n24575 ;
  assign n24550 = n24537 ^ n24108 ;
  assign n24551 = n24538 & n24550 ;
  assign n24552 = n24551 ^ n24108 ;
  assign n24578 = n24577 ^ n24552 ;
  assign n24579 = n24578 ^ n23194 ;
  assign n24546 = n24539 ^ n24512 ;
  assign n24547 = ~n24513 & n24546 ;
  assign n24548 = n24547 ^ n22529 ;
  assign n24549 = n24548 ^ n22571 ;
  assign n24580 = n24579 ^ n24549 ;
  assign n24582 = n24580 ^ x228 ;
  assign n24581 = n24580 ^ n24540 ;
  assign n24583 = n24582 ^ n24581 ;
  assign n24584 = n24545 & ~n24583 ;
  assign n24585 = n24584 ^ n24582 ;
  assign n24611 = n24577 ^ n24114 ;
  assign n24612 = n24578 & ~n24611 ;
  assign n24613 = n24612 ^ n24114 ;
  assign n24609 = ~n24575 & n24576 ;
  assign n24591 = n24561 ^ n24555 ;
  assign n24592 = n24560 & ~n24591 ;
  assign n24593 = n24592 ^ n24555 ;
  assign n24590 = n23967 ^ n23966 ;
  assign n24594 = n24593 ^ n24590 ;
  assign n24595 = n24594 ^ n23842 ;
  assign n24596 = n24595 ^ n23843 ;
  assign n24598 = n24596 ^ n23247 ;
  assign n24597 = n24596 ^ n24563 ;
  assign n24599 = n24598 ^ n24597 ;
  assign n24600 = ~n24568 & n24599 ;
  assign n24601 = n24600 ^ n24598 ;
  assign n24602 = n24601 ^ n22802 ;
  assign n24604 = n24602 ^ x158 ;
  assign n24603 = n24602 ^ n24569 ;
  assign n24605 = n24604 ^ n24603 ;
  assign n24606 = ~n24574 & n24605 ;
  assign n24607 = n24606 ^ n24604 ;
  assign n24608 = n24607 ^ x157 ;
  assign n24610 = n24609 ^ n24608 ;
  assign n24614 = n24613 ^ n24610 ;
  assign n24615 = n24614 ^ n23189 ;
  assign n24586 = n24579 ^ n24548 ;
  assign n24587 = n24549 & ~n24586 ;
  assign n24588 = n24587 ^ n22571 ;
  assign n24589 = n24588 ^ n22612 ;
  assign n24616 = n24615 ^ n24589 ;
  assign n24618 = n24616 ^ x227 ;
  assign n24617 = n24616 ^ n24580 ;
  assign n24619 = n24618 ^ n24617 ;
  assign n24620 = ~n24585 & n24619 ;
  assign n24621 = n24620 ^ n24618 ;
  assign n24649 = n24608 & ~n24609 ;
  assign n24639 = n23969 ^ n23968 ;
  assign n24635 = n23865 ^ n23842 ;
  assign n24634 = n24593 ^ n23865 ;
  assign n24636 = n24635 ^ n24634 ;
  assign n24637 = ~n24594 & ~n24636 ;
  assign n24638 = n24637 ^ n24635 ;
  assign n24640 = n24639 ^ n24638 ;
  assign n24641 = n24640 ^ n23866 ;
  assign n24630 = n24596 ^ n22802 ;
  assign n24631 = n24601 & n24630 ;
  assign n24632 = n24631 ^ n22802 ;
  assign n24633 = n24632 ^ n22847 ;
  assign n24642 = n24641 ^ n24633 ;
  assign n24644 = n24642 ^ x157 ;
  assign n24643 = n24642 ^ n24602 ;
  assign n24645 = n24644 ^ n24643 ;
  assign n24646 = ~n24607 & n24645 ;
  assign n24647 = n24646 ^ n24644 ;
  assign n24648 = n24647 ^ x156 ;
  assign n24650 = n24649 ^ n24648 ;
  assign n24627 = n24613 ^ n24120 ;
  assign n24628 = ~n24614 & ~n24627 ;
  assign n24629 = n24628 ^ n24120 ;
  assign n24651 = n24650 ^ n24629 ;
  assign n24652 = n24651 ^ n24034 ;
  assign n24623 = n24615 ^ n24588 ;
  assign n24624 = ~n24589 & n24623 ;
  assign n24625 = n24624 ^ n22612 ;
  assign n24626 = n24625 ^ n22653 ;
  assign n24653 = n24652 ^ n24626 ;
  assign n24655 = n24653 ^ x226 ;
  assign n24654 = n24653 ^ n24616 ;
  assign n24656 = n24655 ^ n24654 ;
  assign n24657 = ~n24621 & n24656 ;
  assign n24658 = n24657 ^ n24655 ;
  assign n24680 = n23972 ^ n23970 ;
  assign n24674 = n23884 ^ n23332 ;
  assign n24676 = n24674 ^ n23865 ;
  assign n24675 = n24674 ^ n24639 ;
  assign n24677 = n24676 ^ n24675 ;
  assign n24678 = ~n24638 & ~n24677 ;
  assign n24679 = n24678 ^ n24676 ;
  assign n24681 = n24680 ^ n24679 ;
  assign n24682 = n24681 ^ n23884 ;
  assign n24669 = n24641 ^ n24632 ;
  assign n24670 = n24641 ^ n22847 ;
  assign n24671 = ~n24669 & ~n24670 ;
  assign n24672 = n24671 ^ n22847 ;
  assign n24673 = n24672 ^ n22882 ;
  assign n24683 = n24682 ^ n24673 ;
  assign n24685 = n24683 ^ x156 ;
  assign n24684 = n24683 ^ n24642 ;
  assign n24686 = n24685 ^ n24684 ;
  assign n24687 = ~n24647 & n24686 ;
  assign n24688 = n24687 ^ n24685 ;
  assign n24689 = n24688 ^ x155 ;
  assign n24668 = ~n24648 & ~n24649 ;
  assign n24690 = n24689 ^ n24668 ;
  assign n24665 = n24650 ^ n24126 ;
  assign n24666 = n24651 & n24665 ;
  assign n24667 = n24666 ^ n24126 ;
  assign n24691 = n24690 ^ n24667 ;
  assign n24692 = n24691 ^ n23185 ;
  assign n24661 = n24652 ^ n24625 ;
  assign n24662 = ~n24626 & ~n24661 ;
  assign n24663 = n24662 ^ n22653 ;
  assign n24664 = n24663 ^ n22694 ;
  assign n24693 = n24692 ^ n24664 ;
  assign n24695 = n24693 ^ x225 ;
  assign n24694 = n24693 ^ n24653 ;
  assign n24696 = n24695 ^ n24694 ;
  assign n24697 = ~n24658 & n24696 ;
  assign n24698 = n24697 ^ n24695 ;
  assign n24716 = n24680 ^ n24674 ;
  assign n24717 = n24679 & ~n24716 ;
  assign n24715 = n24674 ^ n23903 ;
  assign n24718 = n24717 ^ n24715 ;
  assign n24714 = n23974 ^ n23973 ;
  assign n24719 = n24718 ^ n24714 ;
  assign n24720 = n24719 ^ n23904 ;
  assign n24709 = n24682 ^ n24672 ;
  assign n24710 = n24682 ^ n22882 ;
  assign n24711 = ~n24709 & n24710 ;
  assign n24712 = n24711 ^ n22882 ;
  assign n24713 = n24712 ^ n22920 ;
  assign n24721 = n24720 ^ n24713 ;
  assign n24723 = n24721 ^ x155 ;
  assign n24722 = n24721 ^ n24683 ;
  assign n24724 = n24723 ^ n24722 ;
  assign n24725 = ~n24688 & n24724 ;
  assign n24726 = n24725 ^ n24723 ;
  assign n24727 = n24726 ^ x154 ;
  assign n24708 = ~n24668 & n24689 ;
  assign n24728 = n24727 ^ n24708 ;
  assign n24705 = n24690 ^ n24089 ;
  assign n24706 = ~n24691 & ~n24705 ;
  assign n24707 = n24706 ^ n24089 ;
  assign n24729 = n24728 ^ n24707 ;
  assign n24730 = n24729 ^ n23136 ;
  assign n24701 = n24692 ^ n24663 ;
  assign n24702 = n24664 & ~n24701 ;
  assign n24703 = n24702 ^ n22694 ;
  assign n24704 = n24703 ^ n22735 ;
  assign n24731 = n24730 ^ n24704 ;
  assign n24733 = n24731 ^ x224 ;
  assign n24732 = n24731 ^ n24693 ;
  assign n24734 = n24733 ^ n24732 ;
  assign n24735 = ~n24698 & n24734 ;
  assign n24736 = n24735 ^ n24733 ;
  assign n24766 = n24728 ^ n24136 ;
  assign n24767 = n24729 & ~n24766 ;
  assign n24768 = n24767 ^ n24136 ;
  assign n24755 = n23976 ^ n23975 ;
  assign n24749 = n23922 ^ n23356 ;
  assign n24750 = n24749 ^ n23903 ;
  assign n24751 = n24750 ^ n24714 ;
  assign n24752 = n24751 ^ n24749 ;
  assign n24753 = ~n24718 & n24752 ;
  assign n24754 = n24753 ^ n24750 ;
  assign n24756 = n24755 ^ n24754 ;
  assign n24757 = n24756 ^ n23922 ;
  assign n24744 = n24720 ^ n24712 ;
  assign n24745 = n24720 ^ n22920 ;
  assign n24746 = ~n24744 & ~n24745 ;
  assign n24747 = n24746 ^ n22920 ;
  assign n24748 = n24747 ^ n22967 ;
  assign n24758 = n24757 ^ n24748 ;
  assign n24760 = n24758 ^ x154 ;
  assign n24759 = n24758 ^ n24721 ;
  assign n24761 = n24760 ^ n24759 ;
  assign n24762 = n24726 & ~n24761 ;
  assign n24763 = n24762 ^ n24760 ;
  assign n24764 = n24763 ^ x153 ;
  assign n24743 = n24708 & ~n24727 ;
  assign n24765 = n24764 ^ n24743 ;
  assign n24769 = n24768 ^ n24765 ;
  assign n24770 = n24769 ^ n24047 ;
  assign n24739 = n24730 ^ n24703 ;
  assign n24740 = n24704 & ~n24739 ;
  assign n24741 = n24740 ^ n22735 ;
  assign n24742 = n24741 ^ n22776 ;
  assign n24771 = n24770 ^ n24742 ;
  assign n24773 = n24771 ^ x239 ;
  assign n24772 = n24771 ^ n24731 ;
  assign n24774 = n24773 ^ n24772 ;
  assign n24775 = ~n24736 & n24774 ;
  assign n24776 = n24775 ^ n24773 ;
  assign n24800 = n24758 ^ n24743 ;
  assign n24803 = ~n24763 & ~n24800 ;
  assign n24799 = n24763 ^ n24758 ;
  assign n24801 = n24800 ^ n24799 ;
  assign n24802 = x153 & ~n24801 ;
  assign n24804 = n24803 ^ n24802 ;
  assign n24793 = n24755 ^ n24749 ;
  assign n24794 = n24754 & ~n24793 ;
  assign n24790 = n24010 ^ n23977 ;
  assign n24791 = n24790 ^ n23978 ;
  assign n24792 = n24791 ^ n24755 ;
  assign n24795 = n24794 ^ n24792 ;
  assign n24796 = n24795 ^ n24012 ;
  assign n24789 = n22967 ^ x152 ;
  assign n24797 = n24796 ^ n24789 ;
  assign n24786 = n24757 ^ n24747 ;
  assign n24787 = n24757 ^ n22967 ;
  assign n24788 = ~n24786 & ~n24787 ;
  assign n24798 = n24797 ^ n24788 ;
  assign n24805 = n24804 ^ n24798 ;
  assign n24783 = n24768 ^ n24142 ;
  assign n24784 = n24769 & n24783 ;
  assign n24785 = n24784 ^ n24142 ;
  assign n24806 = n24805 ^ n24785 ;
  assign n24807 = n24806 ^ n24051 ;
  assign n24779 = n24770 ^ n24741 ;
  assign n24780 = ~n24742 & n24779 ;
  assign n24781 = n24780 ^ n22776 ;
  assign n24782 = n24781 ^ n22817 ;
  assign n24808 = n24807 ^ n24782 ;
  assign n24810 = n24808 ^ x238 ;
  assign n24809 = n24808 ^ n24771 ;
  assign n24811 = n24810 ^ n24809 ;
  assign n24812 = ~n24776 & n24811 ;
  assign n24813 = n24812 ^ n24810 ;
  assign n24820 = n24805 ^ n24148 ;
  assign n24821 = n24806 & n24820 ;
  assign n24822 = n24821 ^ n24148 ;
  assign n24823 = n24822 ^ n24397 ;
  assign n24824 = n24823 ^ n24054 ;
  assign n24816 = n24807 ^ n24781 ;
  assign n24817 = n24782 & ~n24816 ;
  assign n24818 = n24817 ^ n22817 ;
  assign n24819 = n24818 ^ n22858 ;
  assign n24825 = n24824 ^ n24819 ;
  assign n24827 = n24825 ^ x237 ;
  assign n24826 = n24825 ^ n24808 ;
  assign n24828 = n24827 ^ n24826 ;
  assign n24829 = n24813 & ~n24828 ;
  assign n24830 = n24829 ^ n24827 ;
  assign n24847 = n24825 ^ x236 ;
  assign n24848 = ~n24830 & n24847 ;
  assign n24849 = n24848 ^ x236 ;
  assign n24842 = n24399 ^ n24397 ;
  assign n24837 = n24160 ^ n24154 ;
  assign n24838 = n24837 ^ n24160 ;
  assign n24839 = n24838 ^ n24822 ;
  assign n24840 = n24823 & ~n24839 ;
  assign n24841 = n24840 ^ n24837 ;
  assign n24843 = n24842 ^ n24841 ;
  assign n24844 = n24843 ^ n24160 ;
  assign n24845 = n24844 ^ n24063 ;
  assign n24833 = n24824 ^ n24818 ;
  assign n24834 = ~n24819 & ~n24833 ;
  assign n24835 = n24834 ^ n22858 ;
  assign n24836 = n24835 ^ n22897 ;
  assign n24846 = n24845 ^ n24836 ;
  assign n24850 = n24849 ^ n24846 ;
  assign n24863 = n24401 ^ n24400 ;
  assign n24859 = n24166 ^ n24160 ;
  assign n24858 = n24842 ^ n24166 ;
  assign n24860 = n24859 ^ n24858 ;
  assign n24861 = n24841 & n24860 ;
  assign n24862 = n24861 ^ n24859 ;
  assign n24864 = n24863 ^ n24862 ;
  assign n24865 = n24864 ^ n24166 ;
  assign n24866 = n24865 ^ n24071 ;
  assign n24853 = n24845 ^ n22897 ;
  assign n24854 = n24845 ^ n24835 ;
  assign n24855 = n24853 & n24854 ;
  assign n24856 = n24855 ^ n22897 ;
  assign n24857 = n24856 ^ n22937 ;
  assign n24867 = n24866 ^ n24857 ;
  assign n24868 = n24867 ^ x235 ;
  assign n24869 = n24868 ^ n24849 ;
  assign n24870 = n24869 ^ n24867 ;
  assign n24871 = ~n24850 & n24870 ;
  assign n24872 = n24871 ^ n24868 ;
  assign n24882 = n24863 ^ n24166 ;
  assign n24883 = n24862 & ~n24882 ;
  assign n24881 = n24166 ^ n24086 ;
  assign n24884 = n24883 ^ n24881 ;
  assign n24880 = n24403 ^ n24402 ;
  assign n24885 = n24884 ^ n24880 ;
  assign n24886 = n24885 ^ n24086 ;
  assign n24887 = n24886 ^ n24079 ;
  assign n24875 = n24866 ^ n22937 ;
  assign n24876 = n24866 ^ n24856 ;
  assign n24877 = n24875 & n24876 ;
  assign n24878 = n24877 ^ n22937 ;
  assign n24879 = n24878 ^ n22979 ;
  assign n24888 = n24887 ^ n24879 ;
  assign n24890 = n24888 ^ x234 ;
  assign n24889 = n24888 ^ n24867 ;
  assign n24891 = n24890 ^ n24889 ;
  assign n24892 = n24872 & ~n24891 ;
  assign n24893 = n24892 ^ n24890 ;
  assign n24904 = n24887 ^ n22979 ;
  assign n24905 = n24887 ^ n24878 ;
  assign n24906 = ~n24904 & ~n24905 ;
  assign n24907 = n24906 ^ n22979 ;
  assign n24908 = n24907 ^ n23020 ;
  assign n24898 = n24880 ^ n24086 ;
  assign n24899 = n24884 & ~n24898 ;
  assign n24897 = n24181 ^ n24086 ;
  assign n24900 = n24899 ^ n24897 ;
  assign n24896 = n24405 ^ n24404 ;
  assign n24901 = n24900 ^ n24896 ;
  assign n24902 = n24901 ^ n24181 ;
  assign n24903 = n24902 ^ n24175 ;
  assign n24909 = n24908 ^ n24903 ;
  assign n24911 = n24909 ^ x233 ;
  assign n24910 = n24909 ^ n24888 ;
  assign n24912 = n24911 ^ n24910 ;
  assign n24913 = n24893 & ~n24912 ;
  assign n24914 = n24913 ^ n24911 ;
  assign n24932 = n24909 ^ x232 ;
  assign n24933 = ~n24914 & n24932 ;
  assign n24934 = n24933 ^ x232 ;
  assign n24935 = n24934 ^ x247 ;
  assign n24917 = n24907 ^ n24903 ;
  assign n24920 = n24896 ^ n24181 ;
  assign n24921 = ~n24900 & n24920 ;
  assign n24922 = n24921 ^ n24181 ;
  assign n24918 = n24406 ^ n24396 ;
  assign n24919 = n24918 ^ n24285 ;
  assign n24923 = n24922 ^ n24919 ;
  assign n24924 = n24923 ^ n24285 ;
  assign n24925 = n24924 ^ n24282 ;
  assign n24926 = n24925 ^ n23020 ;
  assign n24927 = n24926 ^ n24903 ;
  assign n24928 = n24927 ^ n24925 ;
  assign n24929 = n24917 & ~n24928 ;
  assign n24930 = n24929 ^ n24926 ;
  assign n24931 = n24930 ^ n23062 ;
  assign n24936 = n24935 ^ n24931 ;
  assign n24622 = n24621 ^ x226 ;
  assign n24659 = n24658 ^ x225 ;
  assign n24660 = ~n24622 & ~n24659 ;
  assign n24699 = n24698 ^ x224 ;
  assign n24700 = ~n24660 & n24699 ;
  assign n24737 = n24736 ^ x239 ;
  assign n24738 = ~n24700 & ~n24737 ;
  assign n24777 = n24776 ^ x238 ;
  assign n24778 = n24738 & ~n24777 ;
  assign n24814 = n24813 ^ x237 ;
  assign n24815 = ~n24778 & ~n24814 ;
  assign n24831 = n24830 ^ x236 ;
  assign n24832 = ~n24815 & ~n24831 ;
  assign n24851 = n24850 ^ x235 ;
  assign n24852 = ~n24832 & n24851 ;
  assign n24873 = n24872 ^ x234 ;
  assign n24874 = n24852 & ~n24873 ;
  assign n24894 = n24893 ^ x233 ;
  assign n24895 = ~n24874 & n24894 ;
  assign n24915 = n24914 ^ x232 ;
  assign n24916 = ~n24895 & n24915 ;
  assign n24937 = n24936 ^ n24916 ;
  assign n24938 = n24937 ^ n23987 ;
  assign n25650 = x327 & ~n24938 ;
  assign n25222 = ~n24916 & n24936 ;
  assign n25047 = n24934 ^ n24931 ;
  assign n25048 = n24935 & n25047 ;
  assign n25049 = n25048 ^ x247 ;
  assign n25220 = n25049 ^ x246 ;
  assign n24961 = n24294 ^ n23062 ;
  assign n24947 = n24922 ^ n24918 ;
  assign n24945 = n24408 ^ n24407 ;
  assign n24948 = n24945 ^ n24285 ;
  assign n24949 = n24948 ^ n24918 ;
  assign n24950 = n24949 ^ n24945 ;
  assign n24951 = ~n24947 & n24950 ;
  assign n24952 = n24951 ^ n24948 ;
  assign n24962 = n24961 ^ n24952 ;
  assign n24960 = n24925 ^ n24294 ;
  assign n24963 = n24962 ^ n24960 ;
  assign n24964 = n24963 ^ n24952 ;
  assign n24965 = n24930 & n24964 ;
  assign n24966 = n24965 ^ n24962 ;
  assign n25046 = n24966 ^ n23121 ;
  assign n25221 = n25220 ^ n25046 ;
  assign n25249 = n25222 ^ n25221 ;
  assign n25246 = n24499 ^ n24466 ;
  assign n25244 = n24440 ^ n24097 ;
  assign n25245 = n24937 & n25244 ;
  assign n25247 = n25246 ^ n25245 ;
  assign n25401 = n25249 ^ n25247 ;
  assign n25402 = n25401 ^ n24469 ;
  assign n25399 = n24937 ^ n24467 ;
  assign n25400 = ~n23986 & n25399 ;
  assign n25403 = n25402 ^ n25400 ;
  assign n25649 = n25403 ^ n23990 ;
  assign n25651 = n25650 ^ n25649 ;
  assign n25404 = n25400 ^ n23990 ;
  assign n25405 = ~n25403 & ~n25404 ;
  assign n25406 = n25405 ^ n23990 ;
  assign n25652 = n25406 ^ n23197 ;
  assign n25223 = ~n25221 & n25222 ;
  assign n25050 = n25049 ^ n25046 ;
  assign n24959 = n24952 ^ n23546 ;
  assign n24967 = n24959 & n24966 ;
  assign n24946 = n24945 ^ n24300 ;
  assign n24953 = ~n24946 & n24952 ;
  assign n24944 = n24320 ^ n24300 ;
  assign n24954 = n24953 ^ n24944 ;
  assign n24943 = n24410 ^ n24409 ;
  assign n24955 = n24954 ^ n24943 ;
  assign n24956 = n24955 ^ n24320 ;
  assign n24957 = n24956 ^ n24317 ;
  assign n24958 = n24957 ^ n23121 ;
  assign n24968 = n24967 ^ n24958 ;
  assign n25051 = n24968 ^ n23256 ;
  assign n25052 = n25051 ^ x246 ;
  assign n25053 = n25052 ^ n25046 ;
  assign n25054 = n25053 ^ n25051 ;
  assign n25055 = ~n25050 & n25054 ;
  assign n25056 = n25055 ^ n25052 ;
  assign n25219 = n25056 ^ x245 ;
  assign n25258 = n25223 ^ n25219 ;
  assign n25248 = n24514 ^ n24498 ;
  assign n25250 = n25249 ^ n25248 ;
  assign n25251 = n25250 ^ n25246 ;
  assign n25252 = n25251 ^ n25248 ;
  assign n25253 = n25247 & ~n25252 ;
  assign n25254 = n25253 ^ n25250 ;
  assign n25407 = n25258 ^ n25254 ;
  assign n25408 = n25407 ^ n24502 ;
  assign n25653 = n25652 ^ n25408 ;
  assign n25654 = n25653 ^ x326 ;
  assign n25655 = n25654 ^ n25649 ;
  assign n25656 = n25655 ^ n25653 ;
  assign n25657 = n25651 & ~n25656 ;
  assign n25658 = n25657 ^ n25654 ;
  assign n25409 = n25408 ^ n25406 ;
  assign n25410 = n25408 ^ n23197 ;
  assign n25411 = ~n25409 & n25410 ;
  assign n25412 = n25411 ^ n23197 ;
  assign n25659 = n25412 ^ n23998 ;
  assign n25224 = n25219 & ~n25223 ;
  assign n24975 = n24943 ^ n24320 ;
  assign n24976 = n24954 & ~n24975 ;
  assign n24974 = n24345 ^ n24320 ;
  assign n24977 = n24976 ^ n24974 ;
  assign n24973 = n24412 ^ n24411 ;
  assign n24978 = n24977 ^ n24973 ;
  assign n24979 = n24978 ^ n24345 ;
  assign n24980 = n24979 ^ n24338 ;
  assign n24969 = n24957 ^ n23256 ;
  assign n24970 = ~n24968 & ~n24969 ;
  assign n24971 = n24970 ^ n23256 ;
  assign n24972 = n24971 ^ n23266 ;
  assign n25057 = n24980 ^ n24972 ;
  assign n25059 = n25057 ^ x245 ;
  assign n25058 = n25057 ^ n25051 ;
  assign n25060 = n25059 ^ n25058 ;
  assign n25061 = ~n25056 & n25060 ;
  assign n25062 = n25061 ^ n25059 ;
  assign n25218 = n25062 ^ x244 ;
  assign n25266 = n25224 ^ n25218 ;
  assign n25255 = n24516 ^ n24108 ;
  assign n25256 = n25255 ^ n24537 ;
  assign n25259 = n25258 ^ n25256 ;
  assign n25257 = n25256 ^ n25248 ;
  assign n25260 = n25259 ^ n25257 ;
  assign n25261 = ~n25254 & n25260 ;
  assign n25262 = n25261 ^ n25257 ;
  assign n25396 = n25266 ^ n25262 ;
  assign n25397 = n25396 ^ n24538 ;
  assign n25660 = n25659 ^ n25397 ;
  assign n25662 = n25660 ^ x325 ;
  assign n25661 = n25660 ^ n25653 ;
  assign n25663 = n25662 ^ n25661 ;
  assign n25664 = n25658 & ~n25663 ;
  assign n25665 = n25664 ^ n25662 ;
  assign n25225 = n25218 & ~n25224 ;
  assign n24987 = n24973 ^ n24345 ;
  assign n24988 = ~n24977 & n24987 ;
  assign n24986 = n24366 ^ n24345 ;
  assign n24989 = n24988 ^ n24986 ;
  assign n24985 = n24414 ^ n24413 ;
  assign n24990 = n24989 ^ n24985 ;
  assign n24991 = n24990 ^ n24366 ;
  assign n24992 = n24991 ^ n24359 ;
  assign n24981 = n24980 ^ n24971 ;
  assign n24982 = ~n24972 & ~n24981 ;
  assign n24983 = n24982 ^ n23266 ;
  assign n24984 = n24983 ^ n23272 ;
  assign n25063 = n24992 ^ n24984 ;
  assign n25065 = n25063 ^ x244 ;
  assign n25064 = n25063 ^ n25057 ;
  assign n25066 = n25065 ^ n25064 ;
  assign n25067 = n25062 & ~n25066 ;
  assign n25068 = n25067 ^ n25065 ;
  assign n25217 = n25068 ^ x243 ;
  assign n25273 = n25225 ^ n25217 ;
  assign n25263 = n24552 ^ n24114 ;
  assign n25264 = n25263 ^ n24577 ;
  assign n25267 = n25266 ^ n25264 ;
  assign n25265 = n25264 ^ n25256 ;
  assign n25268 = n25267 ^ n25265 ;
  assign n25269 = ~n25262 & n25268 ;
  assign n25270 = n25269 ^ n25265 ;
  assign n25417 = n25273 ^ n25270 ;
  assign n25418 = n25417 ^ n24578 ;
  assign n25398 = n25397 ^ n23998 ;
  assign n25413 = n25412 ^ n25397 ;
  assign n25414 = ~n25398 & n25413 ;
  assign n25415 = n25414 ^ n23998 ;
  assign n25416 = n25415 ^ n23194 ;
  assign n25666 = n25418 ^ n25416 ;
  assign n25668 = n25666 ^ x324 ;
  assign n25667 = n25666 ^ n25660 ;
  assign n25669 = n25668 ^ n25667 ;
  assign n25670 = ~n25665 & n25669 ;
  assign n25671 = n25670 ^ n25668 ;
  assign n25833 = n25671 ^ x323 ;
  assign n25226 = ~n25217 & n25225 ;
  assign n24999 = n24985 ^ n24366 ;
  assign n25000 = n24989 & ~n24999 ;
  assign n24998 = n24387 ^ n24366 ;
  assign n25001 = n25000 ^ n24998 ;
  assign n24997 = n24416 ^ n24415 ;
  assign n25002 = n25001 ^ n24997 ;
  assign n25003 = n25002 ^ n24387 ;
  assign n25004 = n25003 ^ n24380 ;
  assign n24993 = n24992 ^ n24983 ;
  assign n24994 = ~n24984 & ~n24993 ;
  assign n24995 = n24994 ^ n23272 ;
  assign n24996 = n24995 ^ n23278 ;
  assign n25069 = n25004 ^ n24996 ;
  assign n25071 = n25069 ^ x243 ;
  assign n25070 = n25069 ^ n25063 ;
  assign n25072 = n25071 ^ n25070 ;
  assign n25073 = ~n25068 & n25072 ;
  assign n25074 = n25073 ^ n25071 ;
  assign n25216 = n25074 ^ x242 ;
  assign n25281 = n25226 ^ n25216 ;
  assign n25271 = n24627 ^ n24610 ;
  assign n25274 = n25273 ^ n25271 ;
  assign n25272 = n25271 ^ n25264 ;
  assign n25275 = n25274 ^ n25272 ;
  assign n25276 = n25270 & n25275 ;
  assign n25277 = n25276 ^ n25272 ;
  assign n25423 = n25281 ^ n25277 ;
  assign n25424 = n25423 ^ n24614 ;
  assign n25419 = n25418 ^ n25415 ;
  assign n25420 = n25416 & ~n25419 ;
  assign n25421 = n25420 ^ n23194 ;
  assign n25422 = n25421 ^ n23189 ;
  assign n25672 = n25424 ^ n25422 ;
  assign n25674 = n25672 ^ x323 ;
  assign n25673 = n25672 ^ n25666 ;
  assign n25675 = n25674 ^ n25673 ;
  assign n25676 = n25671 & ~n25675 ;
  assign n25677 = n25676 ^ n25674 ;
  assign n25834 = n25677 ^ x322 ;
  assign n25835 = n25833 & n25834 ;
  assign n25227 = n25216 & n25226 ;
  assign n25011 = n24997 ^ n24387 ;
  assign n25012 = ~n25001 & n25011 ;
  assign n25010 = n24456 ^ n24387 ;
  assign n25013 = n25012 ^ n25010 ;
  assign n25009 = n24418 ^ n24417 ;
  assign n25014 = n25013 ^ n25009 ;
  assign n25015 = n25014 ^ n24456 ;
  assign n25016 = n25015 ^ n24449 ;
  assign n25005 = n25004 ^ n24995 ;
  assign n25006 = ~n24996 & ~n25005 ;
  assign n25007 = n25006 ^ n23278 ;
  assign n25008 = n25007 ^ n23284 ;
  assign n25075 = n25016 ^ n25008 ;
  assign n25077 = n25075 ^ x242 ;
  assign n25076 = n25075 ^ n25069 ;
  assign n25078 = n25077 ^ n25076 ;
  assign n25079 = n25074 & ~n25078 ;
  assign n25080 = n25079 ^ n25077 ;
  assign n25215 = n25080 ^ x241 ;
  assign n25288 = n25227 ^ n25215 ;
  assign n25278 = n24629 ^ n24126 ;
  assign n25279 = n25278 ^ n24650 ;
  assign n25282 = n25281 ^ n25279 ;
  assign n25280 = n25279 ^ n25271 ;
  assign n25283 = n25282 ^ n25280 ;
  assign n25284 = n25277 & ~n25283 ;
  assign n25285 = n25284 ^ n25280 ;
  assign n25429 = n25288 ^ n25285 ;
  assign n25430 = n25429 ^ n24651 ;
  assign n25425 = n25424 ^ n25421 ;
  assign n25426 = n25422 & ~n25425 ;
  assign n25427 = n25426 ^ n23189 ;
  assign n25428 = n25427 ^ n24034 ;
  assign n25678 = n25430 ^ n25428 ;
  assign n25680 = n25678 ^ x322 ;
  assign n25679 = n25678 ^ n25672 ;
  assign n25681 = n25680 ^ n25679 ;
  assign n25682 = n25677 & ~n25681 ;
  assign n25683 = n25682 ^ n25680 ;
  assign n25836 = n25683 ^ x321 ;
  assign n25837 = n25835 & n25836 ;
  assign n25228 = n25215 & ~n25227 ;
  assign n25017 = n25016 ^ n25007 ;
  assign n25018 = ~n25008 & ~n25017 ;
  assign n25019 = n25018 ^ n23284 ;
  assign n25043 = n25019 ^ n23290 ;
  assign n25023 = n24488 ^ n24456 ;
  assign n25021 = n25009 ^ n24456 ;
  assign n25022 = ~n25013 & n25021 ;
  assign n25024 = n25023 ^ n25022 ;
  assign n25020 = n24420 ^ n24419 ;
  assign n25025 = n25024 ^ n25020 ;
  assign n25026 = n25025 ^ n24488 ;
  assign n25027 = n25026 ^ n23568 ;
  assign n25044 = n25043 ^ n25027 ;
  assign n25082 = n25044 ^ x241 ;
  assign n25081 = n25075 ^ n25044 ;
  assign n25083 = n25082 ^ n25081 ;
  assign n25084 = ~n25080 & n25083 ;
  assign n25085 = n25084 ^ n25082 ;
  assign n25214 = n25085 ^ x240 ;
  assign n25297 = n25228 ^ n25214 ;
  assign n25286 = n24667 ^ n24089 ;
  assign n25287 = n25286 ^ n24690 ;
  assign n25290 = n25287 ^ n25279 ;
  assign n25289 = n25288 ^ n25287 ;
  assign n25291 = n25290 ^ n25289 ;
  assign n25292 = n25285 & ~n25291 ;
  assign n25293 = n25292 ^ n25290 ;
  assign n25435 = n25297 ^ n25293 ;
  assign n25436 = n25435 ^ n24691 ;
  assign n25431 = n25430 ^ n25427 ;
  assign n25432 = ~n25428 & n25431 ;
  assign n25433 = n25432 ^ n24034 ;
  assign n25434 = n25433 ^ n23185 ;
  assign n25684 = n25436 ^ n25434 ;
  assign n25686 = n25684 ^ x321 ;
  assign n25685 = n25684 ^ n25678 ;
  assign n25687 = n25686 ^ n25685 ;
  assign n25688 = n25683 & ~n25687 ;
  assign n25689 = n25688 ^ n25686 ;
  assign n25838 = n25689 ^ x320 ;
  assign n25839 = ~n25837 & n25838 ;
  assign n25229 = n25214 & ~n25228 ;
  assign n25045 = n25044 ^ x240 ;
  assign n25086 = ~n25045 & n25085 ;
  assign n25087 = n25086 ^ x240 ;
  assign n25212 = n25087 ^ x255 ;
  assign n25028 = n25027 ^ n25019 ;
  assign n25031 = n25020 ^ n24488 ;
  assign n25032 = n25024 & n25031 ;
  assign n25033 = n25032 ^ n24488 ;
  assign n25029 = n24422 ^ n24421 ;
  assign n25030 = n25029 ^ n24527 ;
  assign n25034 = n25033 ^ n25030 ;
  assign n25035 = n25034 ^ n24527 ;
  assign n25036 = n25035 ^ n23675 ;
  assign n25037 = n25036 ^ n23290 ;
  assign n25038 = n25037 ^ n25019 ;
  assign n25039 = n25038 ^ n25036 ;
  assign n25040 = ~n25028 & ~n25039 ;
  assign n25041 = n25040 ^ n25037 ;
  assign n25042 = n25041 ^ n23293 ;
  assign n25213 = n25212 ^ n25042 ;
  assign n25304 = n25229 ^ n25213 ;
  assign n25294 = n24707 ^ n24136 ;
  assign n25295 = n25294 ^ n24728 ;
  assign n25298 = n25297 ^ n25295 ;
  assign n25296 = n25295 ^ n25287 ;
  assign n25299 = n25298 ^ n25296 ;
  assign n25300 = n25293 & n25299 ;
  assign n25301 = n25300 ^ n25296 ;
  assign n25441 = n25304 ^ n25301 ;
  assign n25442 = n25441 ^ n24729 ;
  assign n25437 = n25436 ^ n25433 ;
  assign n25438 = n25434 & ~n25437 ;
  assign n25439 = n25438 ^ n23185 ;
  assign n25440 = n25439 ^ n23136 ;
  assign n25690 = n25442 ^ n25440 ;
  assign n25692 = n25690 ^ x320 ;
  assign n25691 = n25690 ^ n25684 ;
  assign n25693 = n25692 ^ n25691 ;
  assign n25694 = ~n25689 & n25693 ;
  assign n25695 = n25694 ^ n25692 ;
  assign n25840 = n25695 ^ x335 ;
  assign n25841 = n25839 & n25840 ;
  assign n25230 = n25213 & ~n25229 ;
  assign n25088 = n25087 ^ n25042 ;
  assign n25097 = n24555 ^ n23293 ;
  assign n25094 = n24424 ^ n24423 ;
  assign n25090 = n25033 ^ n25029 ;
  assign n25091 = n25033 ^ n24527 ;
  assign n25092 = ~n25090 & n25091 ;
  assign n25093 = n25092 ^ n24527 ;
  assign n25095 = n25094 ^ n25093 ;
  assign n25098 = n25097 ^ n25095 ;
  assign n25089 = n25036 ^ n24555 ;
  assign n25096 = n25095 ^ n25089 ;
  assign n25099 = n25098 ^ n25096 ;
  assign n25100 = ~n25041 & ~n25099 ;
  assign n25101 = n25100 ^ n25098 ;
  assign n25102 = n25101 ^ n23300 ;
  assign n25103 = n25102 ^ x255 ;
  assign n25104 = n25103 ^ n25042 ;
  assign n25105 = n25104 ^ n25102 ;
  assign n25106 = ~n25088 & n25105 ;
  assign n25107 = n25106 ^ n25103 ;
  assign n25211 = n25107 ^ x254 ;
  assign n25311 = n25230 ^ n25211 ;
  assign n25302 = n24783 ^ n24765 ;
  assign n25305 = n25304 ^ n25302 ;
  assign n25303 = n25302 ^ n25295 ;
  assign n25306 = n25305 ^ n25303 ;
  assign n25307 = ~n25301 & n25306 ;
  assign n25308 = n25307 ^ n25303 ;
  assign n25447 = n25311 ^ n25308 ;
  assign n25448 = n25447 ^ n24769 ;
  assign n25443 = n25442 ^ n25439 ;
  assign n25444 = ~n25440 & n25443 ;
  assign n25445 = n25444 ^ n23136 ;
  assign n25446 = n25445 ^ n24047 ;
  assign n25696 = n25448 ^ n25446 ;
  assign n25698 = n25696 ^ x335 ;
  assign n25697 = n25696 ^ n25690 ;
  assign n25699 = n25698 ^ n25697 ;
  assign n25700 = ~n25695 & n25699 ;
  assign n25701 = n25700 ^ n25698 ;
  assign n25832 = n25701 ^ x334 ;
  assign n25923 = n25841 ^ n25832 ;
  assign n26144 = n25923 ^ n24439 ;
  assign n26145 = x423 & n26144 ;
  assign n26360 = n26145 ^ x422 ;
  assign n25231 = n25211 & ~n25230 ;
  assign n25118 = n25095 ^ n23822 ;
  assign n25119 = ~n25101 & ~n25118 ;
  assign n25113 = n24426 ^ n24425 ;
  assign n25108 = n24595 ^ n24562 ;
  assign n25109 = n25108 ^ n24595 ;
  assign n25110 = n25109 ^ n25093 ;
  assign n25111 = n25095 & n25110 ;
  assign n25112 = n25111 ^ n25108 ;
  assign n25114 = n25113 ^ n25112 ;
  assign n25115 = n25114 ^ n24595 ;
  assign n25116 = n25115 ^ n23842 ;
  assign n25117 = n25116 ^ n23300 ;
  assign n25120 = n25119 ^ n25117 ;
  assign n25121 = n25120 ^ n23253 ;
  assign n25123 = n25121 ^ x254 ;
  assign n25122 = n25121 ^ n25102 ;
  assign n25124 = n25123 ^ n25122 ;
  assign n25125 = n25107 & ~n25124 ;
  assign n25126 = n25125 ^ n25123 ;
  assign n25210 = n25126 ^ x253 ;
  assign n25318 = n25231 ^ n25210 ;
  assign n25309 = n24785 ^ n24148 ;
  assign n25310 = n25309 ^ n24805 ;
  assign n25313 = n25310 ^ n25302 ;
  assign n25312 = n25311 ^ n25310 ;
  assign n25314 = n25313 ^ n25312 ;
  assign n25315 = n25308 & ~n25314 ;
  assign n25316 = n25315 ^ n25313 ;
  assign n25453 = n25318 ^ n25316 ;
  assign n25454 = n25453 ^ n24806 ;
  assign n25449 = n25448 ^ n25445 ;
  assign n25450 = ~n25446 & ~n25449 ;
  assign n25451 = n25450 ^ n24047 ;
  assign n25452 = n25451 ^ n24051 ;
  assign n25702 = n25454 ^ n25452 ;
  assign n25704 = n25702 ^ x334 ;
  assign n25703 = n25702 ^ n25696 ;
  assign n25705 = n25704 ^ n25703 ;
  assign n25706 = ~n25701 & n25705 ;
  assign n25707 = n25706 ^ n25704 ;
  assign n25843 = n25707 ^ x333 ;
  assign n25842 = n25832 & n25841 ;
  assign n25927 = n25843 ^ n25842 ;
  assign n25924 = n25244 ^ n24937 ;
  assign n25925 = n25923 & n25924 ;
  assign n25928 = n25927 ^ n25925 ;
  assign n26028 = n25928 ^ n25246 ;
  assign n26025 = n25923 ^ n25244 ;
  assign n26026 = n24467 & n26025 ;
  assign n26029 = n26028 ^ n26026 ;
  assign n26143 = n26029 ^ n24095 ;
  assign n26361 = n26360 ^ n26143 ;
  assign n26146 = n26145 ^ n26143 ;
  assign n26027 = n26026 ^ n24095 ;
  assign n26030 = n26027 & n26029 ;
  assign n26031 = n26030 ^ n24095 ;
  assign n26147 = n26031 ^ n24092 ;
  assign n25926 = n25925 ^ n25401 ;
  assign n25929 = ~n25926 & ~n25928 ;
  assign n25930 = n25929 ^ n25401 ;
  assign n25241 = n24397 ^ n24154 ;
  assign n25242 = n25241 ^ n24822 ;
  assign n25319 = n25318 ^ n25242 ;
  assign n25317 = n25310 ^ n25242 ;
  assign n25320 = n25319 ^ n25317 ;
  assign n25321 = ~n25316 & ~n25320 ;
  assign n25322 = n25321 ^ n25317 ;
  assign n25232 = n25210 & n25231 ;
  assign n25136 = n24429 ^ n24427 ;
  assign n25132 = n24640 ^ n24595 ;
  assign n25131 = n25113 ^ n24640 ;
  assign n25133 = n25132 ^ n25131 ;
  assign n25134 = n25112 & ~n25133 ;
  assign n25135 = n25134 ^ n25132 ;
  assign n25137 = n25136 ^ n25135 ;
  assign n25138 = n25137 ^ n24640 ;
  assign n25139 = n25138 ^ n23865 ;
  assign n25127 = n25116 ^ n23253 ;
  assign n25128 = ~n25120 & n25127 ;
  assign n25129 = n25128 ^ n23253 ;
  assign n25130 = n25129 ^ n23320 ;
  assign n25140 = n25139 ^ n25130 ;
  assign n25142 = n25140 ^ x253 ;
  assign n25141 = n25140 ^ n25121 ;
  assign n25143 = n25142 ^ n25141 ;
  assign n25144 = n25126 & ~n25143 ;
  assign n25145 = n25144 ^ n25142 ;
  assign n25209 = n25145 ^ x252 ;
  assign n25240 = n25232 ^ n25209 ;
  assign n25459 = n25322 ^ n25240 ;
  assign n25460 = n25459 ^ n24823 ;
  assign n25455 = n25454 ^ n25451 ;
  assign n25456 = n25452 & n25455 ;
  assign n25457 = n25456 ^ n24051 ;
  assign n25458 = n25457 ^ n24054 ;
  assign n25708 = n25460 ^ n25458 ;
  assign n25710 = n25708 ^ x333 ;
  assign n25709 = n25708 ^ n25702 ;
  assign n25711 = n25710 ^ n25709 ;
  assign n25712 = n25707 & ~n25711 ;
  assign n25713 = n25712 ^ n25710 ;
  assign n25845 = n25713 ^ x332 ;
  assign n25844 = ~n25842 & n25843 ;
  assign n25921 = n25845 ^ n25844 ;
  assign n25931 = n25930 ^ n25921 ;
  assign n26023 = n25931 ^ n25248 ;
  assign n26148 = n26147 ^ n26023 ;
  assign n26149 = n26148 ^ x422 ;
  assign n26150 = n26149 ^ n26143 ;
  assign n26151 = n26150 ^ n26148 ;
  assign n26152 = n26146 & ~n26151 ;
  assign n26153 = n26152 ^ n26149 ;
  assign n26362 = n26153 ^ x421 ;
  assign n26363 = n26361 & n26362 ;
  assign n26024 = n26023 ^ n24092 ;
  assign n26032 = n26031 ^ n26023 ;
  assign n26033 = ~n26024 & n26032 ;
  assign n26034 = n26033 ^ n24092 ;
  assign n26154 = n26034 ^ n24108 ;
  assign n25922 = n25921 ^ n25407 ;
  assign n25932 = ~n25922 & ~n25931 ;
  assign n25933 = n25932 ^ n25407 ;
  assign n25846 = n25844 & n25845 ;
  assign n25243 = n25242 ^ n25240 ;
  assign n25323 = n25243 & ~n25322 ;
  assign n25324 = n25323 ^ n25242 ;
  assign n25465 = n25324 ^ n24843 ;
  assign n25233 = n25209 & ~n25232 ;
  assign n25156 = n24431 ^ n24430 ;
  assign n25152 = n24681 ^ n24640 ;
  assign n25151 = n25136 ^ n24681 ;
  assign n25153 = n25152 ^ n25151 ;
  assign n25154 = ~n25135 & n25153 ;
  assign n25155 = n25154 ^ n25152 ;
  assign n25157 = n25156 ^ n25155 ;
  assign n25158 = n25157 ^ n24681 ;
  assign n25159 = n25158 ^ n24674 ;
  assign n25146 = n25139 ^ n25129 ;
  assign n25147 = n25139 ^ n23320 ;
  assign n25148 = n25146 & ~n25147 ;
  assign n25149 = n25148 ^ n23320 ;
  assign n25150 = n25149 ^ n23332 ;
  assign n25160 = n25159 ^ n25150 ;
  assign n25162 = n25160 ^ x252 ;
  assign n25161 = n25160 ^ n25140 ;
  assign n25163 = n25162 ^ n25161 ;
  assign n25164 = ~n25145 & n25163 ;
  assign n25165 = n25164 ^ n25162 ;
  assign n25208 = n25165 ^ x251 ;
  assign n25238 = n25233 ^ n25208 ;
  assign n25466 = n25465 ^ n25238 ;
  assign n25467 = n25466 ^ n24844 ;
  assign n25461 = n25460 ^ n25457 ;
  assign n25462 = n25458 & n25461 ;
  assign n25463 = n25462 ^ n24054 ;
  assign n25464 = n25463 ^ n24063 ;
  assign n25714 = n25467 ^ n25464 ;
  assign n25716 = n25714 ^ x332 ;
  assign n25715 = n25714 ^ n25708 ;
  assign n25717 = n25716 ^ n25715 ;
  assign n25718 = n25713 & ~n25717 ;
  assign n25719 = n25718 ^ n25716 ;
  assign n25831 = n25719 ^ x331 ;
  assign n25919 = n25846 ^ n25831 ;
  assign n25934 = n25933 ^ n25919 ;
  assign n26021 = n25934 ^ n25256 ;
  assign n26155 = n26154 ^ n26021 ;
  assign n26157 = n26155 ^ x421 ;
  assign n26156 = n26155 ^ n26148 ;
  assign n26158 = n26157 ^ n26156 ;
  assign n26159 = n26153 & ~n26158 ;
  assign n26160 = n26159 ^ n26157 ;
  assign n26364 = n26160 ^ x420 ;
  assign n26365 = ~n26363 & ~n26364 ;
  assign n25847 = ~n25831 & n25846 ;
  assign n25234 = n25208 & ~n25233 ;
  assign n25176 = n24433 ^ n24432 ;
  assign n25172 = n24719 ^ n24681 ;
  assign n25171 = n25156 ^ n24719 ;
  assign n25173 = n25172 ^ n25171 ;
  assign n25174 = ~n25155 & ~n25173 ;
  assign n25175 = n25174 ^ n25172 ;
  assign n25177 = n25176 ^ n25175 ;
  assign n25178 = n25177 ^ n24719 ;
  assign n25179 = n25178 ^ n23903 ;
  assign n25166 = n25159 ^ n25149 ;
  assign n25167 = n25159 ^ n23332 ;
  assign n25168 = ~n25166 & n25167 ;
  assign n25169 = n25168 ^ n23332 ;
  assign n25170 = n25169 ^ n23344 ;
  assign n25180 = n25179 ^ n25170 ;
  assign n25182 = n25180 ^ x251 ;
  assign n25181 = n25180 ^ n25160 ;
  assign n25183 = n25182 ^ n25181 ;
  assign n25184 = n25165 & ~n25183 ;
  assign n25185 = n25184 ^ n25182 ;
  assign n25207 = n25185 ^ x250 ;
  assign n25329 = n25234 ^ n25207 ;
  assign n25239 = n25238 ^ n24843 ;
  assign n25325 = n25324 ^ n25238 ;
  assign n25326 = n25239 & n25325 ;
  assign n25327 = n25326 ^ n24843 ;
  assign n25328 = n25327 ^ n24864 ;
  assign n25472 = n25329 ^ n25328 ;
  assign n25473 = n25472 ^ n24865 ;
  assign n25468 = n25467 ^ n25463 ;
  assign n25469 = ~n25464 & n25468 ;
  assign n25470 = n25469 ^ n24063 ;
  assign n25471 = n25470 ^ n24071 ;
  assign n25720 = n25473 ^ n25471 ;
  assign n25722 = n25720 ^ x331 ;
  assign n25721 = n25720 ^ n25714 ;
  assign n25723 = n25722 ^ n25721 ;
  assign n25724 = ~n25719 & n25723 ;
  assign n25725 = n25724 ^ n25722 ;
  assign n25830 = n25725 ^ x330 ;
  assign n25938 = n25847 ^ n25830 ;
  assign n25920 = n25919 ^ n25396 ;
  assign n25935 = ~n25920 & ~n25934 ;
  assign n25936 = n25935 ^ n25396 ;
  assign n25939 = n25938 ^ n25936 ;
  assign n26039 = n25939 ^ n25264 ;
  assign n26022 = n26021 ^ n24108 ;
  assign n26035 = n26034 ^ n26021 ;
  assign n26036 = ~n26022 & ~n26035 ;
  assign n26037 = n26036 ^ n24108 ;
  assign n26038 = n26037 ^ n24114 ;
  assign n26141 = n26039 ^ n26038 ;
  assign n26162 = n26141 ^ x420 ;
  assign n26161 = n26155 ^ n26141 ;
  assign n26163 = n26162 ^ n26161 ;
  assign n26164 = n26160 & ~n26163 ;
  assign n26165 = n26164 ^ n26162 ;
  assign n26366 = n26165 ^ x419 ;
  assign n26367 = n26365 & ~n26366 ;
  assign n25937 = n25936 ^ n25417 ;
  assign n25940 = ~n25937 & n25939 ;
  assign n25941 = n25940 ^ n25417 ;
  assign n25474 = n25473 ^ n25470 ;
  assign n25475 = n25471 & n25474 ;
  assign n25476 = n25475 ^ n24071 ;
  assign n25726 = n25476 ^ n24079 ;
  assign n25330 = n25329 ^ n25327 ;
  assign n25331 = ~n25328 & ~n25330 ;
  assign n25332 = n25331 ^ n24864 ;
  assign n25392 = n25332 ^ n24885 ;
  assign n25235 = ~n25207 & n25234 ;
  assign n25196 = n24435 ^ n24434 ;
  assign n25192 = n24756 ^ n24719 ;
  assign n25191 = n25176 ^ n24756 ;
  assign n25193 = n25192 ^ n25191 ;
  assign n25194 = ~n25175 & ~n25193 ;
  assign n25195 = n25194 ^ n25192 ;
  assign n25197 = n25196 ^ n25195 ;
  assign n25198 = n25197 ^ n24756 ;
  assign n25199 = n25198 ^ n24749 ;
  assign n25186 = n25179 ^ n25169 ;
  assign n25187 = n25179 ^ n23344 ;
  assign n25188 = n25186 & ~n25187 ;
  assign n25189 = n25188 ^ n23344 ;
  assign n25190 = n25189 ^ n23356 ;
  assign n25200 = n25199 ^ n25190 ;
  assign n25202 = n25200 ^ x250 ;
  assign n25201 = n25200 ^ n25180 ;
  assign n25203 = n25202 ^ n25201 ;
  assign n25204 = ~n25185 & n25203 ;
  assign n25205 = n25204 ^ n25202 ;
  assign n25206 = n25205 ^ x249 ;
  assign n25236 = n25235 ^ n25206 ;
  assign n25393 = n25392 ^ n25236 ;
  assign n25394 = n25393 ^ n24886 ;
  assign n25727 = n25726 ^ n25394 ;
  assign n25729 = n25727 ^ x330 ;
  assign n25728 = n25727 ^ n25720 ;
  assign n25730 = n25729 ^ n25728 ;
  assign n25731 = ~n25725 & n25730 ;
  assign n25732 = n25731 ^ n25729 ;
  assign n25849 = n25732 ^ x329 ;
  assign n25848 = ~n25830 & n25847 ;
  assign n25917 = n25849 ^ n25848 ;
  assign n25942 = n25941 ^ n25917 ;
  assign n26044 = n25942 ^ n25271 ;
  assign n26040 = n26039 ^ n26037 ;
  assign n26041 = n26038 & ~n26040 ;
  assign n26042 = n26041 ^ n24114 ;
  assign n26043 = n26042 ^ n24120 ;
  assign n26168 = n26044 ^ n26043 ;
  assign n26142 = n26141 ^ x419 ;
  assign n26166 = ~n26142 & n26165 ;
  assign n26167 = n26166 ^ x419 ;
  assign n26169 = n26168 ^ n26167 ;
  assign n26368 = n26169 ^ x418 ;
  assign n26369 = n26367 & n26368 ;
  assign n25918 = n25917 ^ n25423 ;
  assign n25943 = n25918 & n25942 ;
  assign n25944 = n25943 ^ n25423 ;
  assign n25395 = n25394 ^ n24079 ;
  assign n25477 = n25476 ^ n25394 ;
  assign n25478 = ~n25395 & n25477 ;
  assign n25479 = n25478 ^ n24079 ;
  assign n25646 = n25479 ^ n24175 ;
  assign n25354 = n25235 ^ n25200 ;
  assign n25355 = n25205 & ~n25354 ;
  assign n25352 = n25235 ^ n25205 ;
  assign n25353 = x249 & ~n25352 ;
  assign n25356 = n25355 ^ n25353 ;
  assign n25344 = n25196 ^ n24756 ;
  assign n25345 = ~n25195 & n25344 ;
  assign n25341 = n24795 ^ n24437 ;
  assign n25342 = n25341 ^ n24436 ;
  assign n25343 = n25342 ^ n25196 ;
  assign n25346 = n25345 ^ n25343 ;
  assign n25347 = n25346 ^ n24795 ;
  assign n25348 = n25347 ^ n24010 ;
  assign n25349 = n25348 ^ n23367 ;
  assign n25340 = n23356 ^ x248 ;
  assign n25350 = n25349 ^ n25340 ;
  assign n25337 = n25199 ^ n25189 ;
  assign n25338 = n25199 ^ n23356 ;
  assign n25339 = ~n25337 & n25338 ;
  assign n25351 = n25350 ^ n25339 ;
  assign n25357 = n25356 ^ n25351 ;
  assign n25237 = n25236 ^ n24885 ;
  assign n25333 = n25332 ^ n25236 ;
  assign n25334 = n25237 & ~n25333 ;
  assign n25335 = n25334 ^ n24885 ;
  assign n25336 = n25335 ^ n24901 ;
  assign n25480 = n25357 ^ n25336 ;
  assign n25481 = n25480 ^ n24902 ;
  assign n25647 = n25646 ^ n25481 ;
  assign n25734 = n25647 ^ x329 ;
  assign n25733 = n25727 ^ n25647 ;
  assign n25735 = n25734 ^ n25733 ;
  assign n25736 = ~n25732 & n25735 ;
  assign n25737 = n25736 ^ n25734 ;
  assign n25851 = n25737 ^ x328 ;
  assign n25850 = ~n25848 & n25849 ;
  assign n25915 = n25851 ^ n25850 ;
  assign n25945 = n25944 ^ n25915 ;
  assign n26049 = n25945 ^ n25279 ;
  assign n26045 = n26044 ^ n26042 ;
  assign n26046 = ~n26043 & ~n26045 ;
  assign n26047 = n26046 ^ n24120 ;
  assign n26048 = n26047 ^ n24126 ;
  assign n26170 = n26049 ^ n26048 ;
  assign n26171 = n26170 ^ x418 ;
  assign n26172 = n26171 ^ n26167 ;
  assign n26173 = n26172 ^ n26170 ;
  assign n26174 = ~n26169 & n26173 ;
  assign n26175 = n26174 ^ n26171 ;
  assign n26370 = n26175 ^ x417 ;
  assign n26371 = ~n26369 & n26370 ;
  assign n25916 = n25915 ^ n25429 ;
  assign n25946 = n25916 & ~n25945 ;
  assign n25947 = n25946 ^ n25429 ;
  assign n25648 = n25647 ^ x328 ;
  assign n25738 = n25648 & ~n25737 ;
  assign n25739 = n25738 ^ x328 ;
  assign n25853 = n25739 ^ x343 ;
  assign n25482 = n25481 ^ n25479 ;
  assign n25358 = n25357 ^ n25335 ;
  assign n25359 = ~n25336 & n25358 ;
  assign n25360 = n25359 ^ n24901 ;
  assign n24941 = n24440 ^ x231 ;
  assign n24942 = n24941 ^ n24923 ;
  assign n25483 = n25360 ^ n24942 ;
  assign n25484 = n25483 ^ n24924 ;
  assign n25485 = n25484 ^ n24175 ;
  assign n25486 = n25485 ^ n25479 ;
  assign n25487 = n25486 ^ n25484 ;
  assign n25488 = n25482 & n25487 ;
  assign n25489 = n25488 ^ n25485 ;
  assign n25740 = n25489 ^ n24282 ;
  assign n25854 = n25853 ^ n25740 ;
  assign n25852 = ~n25850 & ~n25851 ;
  assign n25913 = n25854 ^ n25852 ;
  assign n25948 = n25947 ^ n25913 ;
  assign n26054 = n25948 ^ n25287 ;
  assign n26050 = n26049 ^ n26047 ;
  assign n26051 = ~n26048 & ~n26050 ;
  assign n26052 = n26051 ^ n24126 ;
  assign n26053 = n26052 ^ n24089 ;
  assign n26176 = n26054 ^ n26053 ;
  assign n26178 = n26176 ^ x417 ;
  assign n26177 = n26176 ^ n26170 ;
  assign n26179 = n26178 ^ n26177 ;
  assign n26180 = n26175 & ~n26179 ;
  assign n26181 = n26180 ^ n26178 ;
  assign n26372 = n26181 ^ x416 ;
  assign n26373 = n26371 & n26372 ;
  assign n25914 = n25913 ^ n25435 ;
  assign n25949 = ~n25914 & ~n25948 ;
  assign n25950 = n25949 ^ n25435 ;
  assign n25741 = n25740 ^ n25739 ;
  assign n25365 = n24952 ^ n24300 ;
  assign n25361 = n25360 ^ n24941 ;
  assign n25362 = n24942 & n25361 ;
  assign n25363 = n25362 ^ n24923 ;
  assign n24940 = n24473 ^ x230 ;
  assign n25364 = n25363 ^ n24940 ;
  assign n25490 = n25365 ^ n25364 ;
  assign n25491 = n25490 ^ n24952 ;
  assign n25493 = n25491 ^ n24282 ;
  assign n25492 = n25491 ^ n25484 ;
  assign n25494 = n25493 ^ n25492 ;
  assign n25495 = n25489 & n25494 ;
  assign n25496 = n25495 ^ n25493 ;
  assign n25742 = n25496 ^ n24294 ;
  assign n25743 = n25742 ^ x343 ;
  assign n25744 = n25743 ^ n25739 ;
  assign n25745 = n25744 ^ n25742 ;
  assign n25746 = n25741 & n25745 ;
  assign n25747 = n25746 ^ n25743 ;
  assign n25856 = n25747 ^ x342 ;
  assign n25855 = n25852 & n25854 ;
  assign n25911 = n25856 ^ n25855 ;
  assign n25951 = n25950 ^ n25911 ;
  assign n26059 = n25951 ^ n25295 ;
  assign n26055 = n26054 ^ n26052 ;
  assign n26056 = ~n26053 & n26055 ;
  assign n26057 = n26056 ^ n24089 ;
  assign n26058 = n26057 ^ n24136 ;
  assign n26182 = n26059 ^ n26058 ;
  assign n26184 = n26182 ^ x416 ;
  assign n26183 = n26182 ^ n26176 ;
  assign n26185 = n26184 ^ n26183 ;
  assign n26186 = n26181 & ~n26185 ;
  assign n26187 = n26186 ^ n26184 ;
  assign n26374 = n26187 ^ x431 ;
  assign n26375 = ~n26373 & n26374 ;
  assign n25912 = n25911 ^ n25441 ;
  assign n25952 = ~n25912 & n25951 ;
  assign n25953 = n25952 ^ n25441 ;
  assign n25368 = n24509 ^ x229 ;
  assign n25369 = n25368 ^ n25363 ;
  assign n25366 = n25365 ^ n25363 ;
  assign n25367 = n25364 & ~n25366 ;
  assign n25370 = n25369 ^ n25367 ;
  assign n25389 = n25370 ^ n24955 ;
  assign n25390 = n25389 ^ n24956 ;
  assign n25498 = n25390 ^ n24294 ;
  assign n25497 = n25491 ^ n25390 ;
  assign n25499 = n25498 ^ n25497 ;
  assign n25500 = n25496 & ~n25499 ;
  assign n25501 = n25500 ^ n25498 ;
  assign n25748 = n25501 ^ n24317 ;
  assign n25750 = n25748 ^ x342 ;
  assign n25749 = n25748 ^ n25742 ;
  assign n25751 = n25750 ^ n25749 ;
  assign n25752 = n25747 & ~n25751 ;
  assign n25753 = n25752 ^ n25750 ;
  assign n25858 = n25753 ^ x341 ;
  assign n25857 = n25855 & n25856 ;
  assign n25909 = n25858 ^ n25857 ;
  assign n25954 = n25953 ^ n25909 ;
  assign n26064 = n25954 ^ n25302 ;
  assign n26060 = n26059 ^ n26057 ;
  assign n26061 = n26058 & ~n26060 ;
  assign n26062 = n26061 ^ n24136 ;
  assign n26063 = n26062 ^ n24142 ;
  assign n26188 = n26064 ^ n26063 ;
  assign n26190 = n26188 ^ x431 ;
  assign n26189 = n26188 ^ n26182 ;
  assign n26191 = n26190 ^ n26189 ;
  assign n26192 = ~n26187 & n26191 ;
  assign n26193 = n26192 ^ n26190 ;
  assign n26376 = n26193 ^ x430 ;
  assign n26377 = ~n26375 & n26376 ;
  assign n25910 = n25909 ^ n25447 ;
  assign n25955 = n25910 & ~n25954 ;
  assign n25956 = n25955 ^ n25447 ;
  assign n25391 = n25390 ^ n24317 ;
  assign n25502 = n25391 & ~n25501 ;
  assign n25503 = n25502 ^ n24317 ;
  assign n25754 = n25503 ^ n24338 ;
  assign n25376 = n24545 ^ x228 ;
  assign n25372 = n24978 ^ n24955 ;
  assign n25371 = n25368 ^ n24978 ;
  assign n25373 = n25372 ^ n25371 ;
  assign n25374 = n25370 & n25373 ;
  assign n25375 = n25374 ^ n25372 ;
  assign n25386 = n25376 ^ n25375 ;
  assign n25387 = n25386 ^ n24979 ;
  assign n25755 = n25754 ^ n25387 ;
  assign n25757 = n25755 ^ x341 ;
  assign n25756 = n25755 ^ n25748 ;
  assign n25758 = n25757 ^ n25756 ;
  assign n25759 = ~n25753 & n25758 ;
  assign n25760 = n25759 ^ n25757 ;
  assign n25860 = n25760 ^ x340 ;
  assign n25859 = n25857 & ~n25858 ;
  assign n25907 = n25860 ^ n25859 ;
  assign n25957 = n25956 ^ n25907 ;
  assign n26069 = n25957 ^ n25310 ;
  assign n26065 = n26064 ^ n26062 ;
  assign n26066 = n26063 & n26065 ;
  assign n26067 = n26066 ^ n24142 ;
  assign n26068 = n26067 ^ n24148 ;
  assign n26194 = n26069 ^ n26068 ;
  assign n26196 = n26194 ^ x430 ;
  assign n26195 = n26194 ^ n26188 ;
  assign n26197 = n26196 ^ n26195 ;
  assign n26198 = n26193 & ~n26197 ;
  assign n26199 = n26198 ^ n26196 ;
  assign n26378 = n26199 ^ x429 ;
  assign n26379 = n26377 & n26378 ;
  assign n25908 = n25907 ^ n25453 ;
  assign n25958 = n25908 & ~n25957 ;
  assign n25959 = n25958 ^ n25453 ;
  assign n25388 = n25387 ^ n24338 ;
  assign n25504 = n25503 ^ n25387 ;
  assign n25505 = n25388 & n25504 ;
  assign n25506 = n25505 ^ n24338 ;
  assign n25761 = n25506 ^ n24359 ;
  assign n25382 = n24585 ^ x227 ;
  assign n25378 = n24990 ^ n24978 ;
  assign n25377 = n25376 ^ n24990 ;
  assign n25379 = n25378 ^ n25377 ;
  assign n25380 = ~n25375 & n25379 ;
  assign n25381 = n25380 ^ n25378 ;
  assign n25383 = n25382 ^ n25381 ;
  assign n25384 = n25383 ^ n24991 ;
  assign n25762 = n25761 ^ n25384 ;
  assign n25764 = n25762 ^ x340 ;
  assign n25763 = n25762 ^ n25755 ;
  assign n25765 = n25764 ^ n25763 ;
  assign n25766 = ~n25760 & n25765 ;
  assign n25767 = n25766 ^ n25764 ;
  assign n25862 = n25767 ^ x339 ;
  assign n25861 = n25859 & ~n25860 ;
  assign n25905 = n25862 ^ n25861 ;
  assign n25960 = n25959 ^ n25905 ;
  assign n26074 = n25960 ^ n25242 ;
  assign n26070 = n26069 ^ n26067 ;
  assign n26071 = ~n26068 & ~n26070 ;
  assign n26072 = n26071 ^ n24148 ;
  assign n26073 = n26072 ^ n24154 ;
  assign n26200 = n26074 ^ n26073 ;
  assign n26202 = n26200 ^ x429 ;
  assign n26201 = n26200 ^ n26194 ;
  assign n26203 = n26202 ^ n26201 ;
  assign n26204 = n26199 & ~n26203 ;
  assign n26205 = n26204 ^ n26202 ;
  assign n26359 = n26205 ^ x428 ;
  assign n26655 = n26379 ^ n26359 ;
  assign n26559 = n25941 ^ n25423 ;
  assign n26560 = n26559 ^ n25917 ;
  assign n26538 = n25938 ^ n25937 ;
  assign n26496 = n25933 ^ n25396 ;
  assign n26497 = n26496 ^ n25919 ;
  assign n26539 = n26538 ^ n26497 ;
  assign n25538 = n24699 ^ n24660 ;
  assign n25511 = n25382 ^ n24990 ;
  assign n25512 = n25381 & ~n25511 ;
  assign n25513 = n25512 ^ n24990 ;
  assign n25521 = n25513 ^ n25002 ;
  assign n25522 = n25014 ^ n24622 ;
  assign n25523 = n25522 ^ n25014 ;
  assign n25524 = n25523 ^ n25513 ;
  assign n25525 = n25521 & n25524 ;
  assign n25526 = n25525 ^ n25522 ;
  assign n25534 = n25025 ^ n25014 ;
  assign n25527 = n24659 ^ n24622 ;
  assign n25533 = n25527 ^ n25025 ;
  assign n25535 = n25534 ^ n25533 ;
  assign n25536 = n25526 & n25535 ;
  assign n25537 = n25536 ^ n25534 ;
  assign n25539 = n25538 ^ n25537 ;
  assign n25540 = n25539 ^ n25026 ;
  assign n25385 = n25384 ^ n24359 ;
  assign n25507 = n25506 ^ n25384 ;
  assign n25508 = ~n25385 & ~n25507 ;
  assign n25509 = n25508 ^ n24359 ;
  assign n25510 = n25509 ^ n24380 ;
  assign n25514 = n25002 ^ n24622 ;
  assign n25515 = n25514 ^ n25513 ;
  assign n25516 = n25515 ^ n25003 ;
  assign n25517 = n25516 ^ n25509 ;
  assign n25518 = ~n25510 & n25517 ;
  assign n25519 = n25518 ^ n24380 ;
  assign n25520 = n25519 ^ n24449 ;
  assign n25528 = n25527 ^ n25526 ;
  assign n25529 = n25528 ^ n25015 ;
  assign n25530 = n25529 ^ n25519 ;
  assign n25531 = ~n25520 & n25530 ;
  assign n25532 = n25531 ^ n24449 ;
  assign n25541 = n25540 ^ n25532 ;
  assign n25547 = n24737 ^ n24700 ;
  assign n25543 = n25034 ^ n25025 ;
  assign n25542 = n25538 ^ n25034 ;
  assign n25544 = n25543 ^ n25542 ;
  assign n25545 = ~n25537 & ~n25544 ;
  assign n25546 = n25545 ^ n25543 ;
  assign n25548 = n25547 ^ n25546 ;
  assign n25549 = n25548 ^ n25035 ;
  assign n25550 = n25549 ^ n23568 ;
  assign n25551 = n25550 ^ n25532 ;
  assign n25552 = n25551 ^ n25549 ;
  assign n25553 = ~n25541 & n25552 ;
  assign n25554 = n25553 ^ n25550 ;
  assign n25784 = n25554 ^ n23675 ;
  assign n25641 = n25532 ^ n23568 ;
  assign n25642 = n25641 ^ n25540 ;
  assign n25643 = n25642 ^ x336 ;
  assign n25775 = n25529 ^ n25520 ;
  assign n25644 = n25516 ^ n25510 ;
  assign n25645 = n25644 ^ x338 ;
  assign n25769 = n25644 ^ x339 ;
  assign n25768 = n25762 ^ n25644 ;
  assign n25770 = n25769 ^ n25768 ;
  assign n25771 = ~n25767 & n25770 ;
  assign n25772 = n25771 ^ n25769 ;
  assign n25773 = n25645 & ~n25772 ;
  assign n25774 = n25773 ^ x338 ;
  assign n25776 = n25775 ^ n25774 ;
  assign n25778 = n25642 ^ x337 ;
  assign n25777 = n25774 ^ n25642 ;
  assign n25779 = n25778 ^ n25777 ;
  assign n25780 = n25776 & n25779 ;
  assign n25781 = n25780 ^ n25778 ;
  assign n25782 = n25643 & ~n25781 ;
  assign n25783 = n25782 ^ x336 ;
  assign n25785 = n25784 ^ n25783 ;
  assign n25560 = n25095 ^ n24562 ;
  assign n25556 = n25547 ^ n25034 ;
  assign n25557 = n25546 & ~n25556 ;
  assign n25558 = n25557 ^ n25034 ;
  assign n25555 = n24777 ^ n24738 ;
  assign n25559 = n25558 ^ n25555 ;
  assign n25561 = n25560 ^ n25559 ;
  assign n25562 = n25561 ^ n25095 ;
  assign n25564 = n25562 ^ n23675 ;
  assign n25563 = n25562 ^ n25549 ;
  assign n25565 = n25564 ^ n25563 ;
  assign n25566 = n25554 & n25565 ;
  assign n25567 = n25566 ^ n25564 ;
  assign n25786 = n25567 ^ n24555 ;
  assign n25787 = n25786 ^ x351 ;
  assign n25788 = n25787 ^ n25783 ;
  assign n25789 = n25788 ^ n25786 ;
  assign n25790 = ~n25785 & n25789 ;
  assign n25791 = n25790 ^ n25787 ;
  assign n25568 = n24814 ^ n24778 ;
  assign n25569 = n25568 ^ n25560 ;
  assign n25570 = n25569 ^ n25558 ;
  assign n25571 = n25570 ^ n25568 ;
  assign n25572 = ~n25559 & ~n25571 ;
  assign n25573 = n25572 ^ n25569 ;
  assign n25574 = n25573 ^ n25114 ;
  assign n25575 = n25574 ^ n25115 ;
  assign n25577 = n25575 ^ n24555 ;
  assign n25576 = n25575 ^ n25562 ;
  assign n25578 = n25577 ^ n25576 ;
  assign n25579 = n25567 & ~n25578 ;
  assign n25580 = n25579 ^ n25577 ;
  assign n25792 = n25580 ^ n23842 ;
  assign n25794 = n25792 ^ x350 ;
  assign n25793 = n25792 ^ n25786 ;
  assign n25795 = n25794 ^ n25793 ;
  assign n25796 = ~n25791 & n25795 ;
  assign n25797 = n25796 ^ n25794 ;
  assign n25581 = n25573 ^ n24594 ;
  assign n25582 = ~n25580 & ~n25581 ;
  assign n25583 = n25582 ^ n23842 ;
  assign n25798 = n25583 ^ n23865 ;
  assign n25589 = n24831 ^ n24815 ;
  assign n25585 = n25137 ^ n25114 ;
  assign n25584 = n25568 ^ n25137 ;
  assign n25586 = n25585 ^ n25584 ;
  assign n25587 = n25573 & ~n25586 ;
  assign n25588 = n25587 ^ n25585 ;
  assign n25590 = n25589 ^ n25588 ;
  assign n25591 = n25590 ^ n25138 ;
  assign n25799 = n25798 ^ n25591 ;
  assign n25801 = n25799 ^ x349 ;
  assign n25800 = n25799 ^ n25792 ;
  assign n25802 = n25801 ^ n25800 ;
  assign n25803 = ~n25797 & n25802 ;
  assign n25804 = n25803 ^ n25801 ;
  assign n25592 = n25591 ^ n25583 ;
  assign n25593 = n25591 ^ n23865 ;
  assign n25594 = n25592 & n25593 ;
  assign n25595 = n25594 ^ n23865 ;
  assign n25805 = n25595 ^ n24674 ;
  assign n25601 = n24851 ^ n24832 ;
  assign n25597 = n25157 ^ n25137 ;
  assign n25596 = n25589 ^ n25157 ;
  assign n25598 = n25597 ^ n25596 ;
  assign n25599 = ~n25588 & ~n25598 ;
  assign n25600 = n25599 ^ n25597 ;
  assign n25602 = n25601 ^ n25600 ;
  assign n25603 = n25602 ^ n25158 ;
  assign n25806 = n25805 ^ n25603 ;
  assign n25808 = n25806 ^ x348 ;
  assign n25807 = n25806 ^ n25799 ;
  assign n25809 = n25808 ^ n25807 ;
  assign n25810 = ~n25804 & n25809 ;
  assign n25811 = n25810 ^ n25808 ;
  assign n25604 = n25603 ^ n25595 ;
  assign n25605 = n25603 ^ n24674 ;
  assign n25606 = ~n25604 & n25605 ;
  assign n25607 = n25606 ^ n24674 ;
  assign n25812 = n25607 ^ n23903 ;
  assign n25613 = n24873 ^ n24852 ;
  assign n25609 = n25177 ^ n25157 ;
  assign n25608 = n25601 ^ n25177 ;
  assign n25610 = n25609 ^ n25608 ;
  assign n25611 = n25600 & ~n25610 ;
  assign n25612 = n25611 ^ n25609 ;
  assign n25614 = n25613 ^ n25612 ;
  assign n25615 = n25614 ^ n25178 ;
  assign n25813 = n25812 ^ n25615 ;
  assign n25815 = n25813 ^ x347 ;
  assign n25814 = n25813 ^ n25806 ;
  assign n25816 = n25815 ^ n25814 ;
  assign n25817 = n25811 & ~n25816 ;
  assign n25818 = n25817 ^ n25815 ;
  assign n25616 = n25615 ^ n25607 ;
  assign n25617 = n25615 ^ n23903 ;
  assign n25618 = n25616 & n25617 ;
  assign n25619 = n25618 ^ n23903 ;
  assign n25819 = n25619 ^ n24749 ;
  assign n25625 = n24894 ^ n24874 ;
  assign n25621 = n25197 ^ n25177 ;
  assign n25620 = n25613 ^ n25197 ;
  assign n25622 = n25621 ^ n25620 ;
  assign n25623 = ~n25612 & n25622 ;
  assign n25624 = n25623 ^ n25621 ;
  assign n25626 = n25625 ^ n25624 ;
  assign n25627 = n25626 ^ n25198 ;
  assign n25820 = n25819 ^ n25627 ;
  assign n25822 = n25820 ^ x346 ;
  assign n25821 = n25820 ^ n25813 ;
  assign n25823 = n25822 ^ n25821 ;
  assign n25824 = n25818 & ~n25823 ;
  assign n25825 = n25824 ^ n25822 ;
  assign n25886 = n25825 ^ x345 ;
  assign n25827 = n25783 ^ x351 ;
  assign n25828 = n25827 ^ n25784 ;
  assign n25829 = n25781 ^ x336 ;
  assign n25863 = n25861 & ~n25862 ;
  assign n25864 = n25772 ^ x338 ;
  assign n25865 = n25863 & ~n25864 ;
  assign n25866 = n25776 ^ x337 ;
  assign n25867 = ~n25865 & ~n25866 ;
  assign n25868 = ~n25829 & ~n25867 ;
  assign n25869 = n25828 & ~n25868 ;
  assign n25870 = n25791 ^ x350 ;
  assign n25871 = ~n25869 & ~n25870 ;
  assign n25872 = n25797 ^ x349 ;
  assign n25873 = n25871 & ~n25872 ;
  assign n25874 = n25804 ^ x348 ;
  assign n25875 = n25873 & ~n25874 ;
  assign n25876 = n25811 ^ x347 ;
  assign n25877 = n25875 & n25876 ;
  assign n25878 = n25818 ^ x346 ;
  assign n25879 = n25877 & n25878 ;
  assign n25887 = n25886 ^ n25879 ;
  assign n25888 = n25887 ^ n25515 ;
  assign n25889 = n25878 ^ n25877 ;
  assign n25890 = n25889 ^ n25383 ;
  assign n25891 = n25876 ^ n25875 ;
  assign n25892 = n25891 ^ n25386 ;
  assign n25893 = n25874 ^ n25873 ;
  assign n25894 = n25893 ^ n25389 ;
  assign n25895 = n25872 ^ n25871 ;
  assign n25896 = n25895 ^ n25490 ;
  assign n25897 = n25870 ^ n25869 ;
  assign n25898 = n25897 ^ n25483 ;
  assign n25899 = n25867 ^ n25829 ;
  assign n25900 = n25899 ^ n25393 ;
  assign n25901 = n25866 ^ n25865 ;
  assign n25902 = n25901 ^ n25472 ;
  assign n25903 = n25864 ^ n25863 ;
  assign n25904 = n25903 ^ n25466 ;
  assign n25906 = n25905 ^ n25459 ;
  assign n25961 = n25906 & ~n25960 ;
  assign n25962 = n25961 ^ n25459 ;
  assign n25963 = n25962 ^ n25903 ;
  assign n25964 = ~n25904 & ~n25963 ;
  assign n25965 = n25964 ^ n25466 ;
  assign n25966 = n25965 ^ n25901 ;
  assign n25967 = ~n25902 & n25966 ;
  assign n25968 = n25967 ^ n25472 ;
  assign n25969 = n25968 ^ n25899 ;
  assign n25970 = n25900 & ~n25969 ;
  assign n25971 = n25970 ^ n25393 ;
  assign n25972 = n25971 ^ n25480 ;
  assign n25973 = n25868 ^ n25828 ;
  assign n25974 = n25973 ^ n25971 ;
  assign n25975 = n25972 & ~n25974 ;
  assign n25976 = n25975 ^ n25480 ;
  assign n25977 = n25976 ^ n25897 ;
  assign n25978 = ~n25898 & ~n25977 ;
  assign n25979 = n25978 ^ n25483 ;
  assign n25980 = n25979 ^ n25895 ;
  assign n25981 = n25896 & ~n25980 ;
  assign n25982 = n25981 ^ n25490 ;
  assign n25983 = n25982 ^ n25893 ;
  assign n25984 = ~n25894 & ~n25983 ;
  assign n25985 = n25984 ^ n25389 ;
  assign n25986 = n25985 ^ n25891 ;
  assign n25987 = ~n25892 & ~n25986 ;
  assign n25988 = n25987 ^ n25386 ;
  assign n25989 = n25988 ^ n25889 ;
  assign n25990 = ~n25890 & n25989 ;
  assign n25991 = n25990 ^ n25383 ;
  assign n25992 = n25991 ^ n25887 ;
  assign n25993 = n25888 & ~n25992 ;
  assign n25994 = n25993 ^ n25515 ;
  assign n25880 = n25879 ^ n25820 ;
  assign n25883 = n25825 & ~n25880 ;
  assign n25826 = n25825 ^ n25820 ;
  assign n25881 = n25880 ^ n25826 ;
  assign n25882 = ~x345 & n25881 ;
  assign n25884 = n25883 ^ n25882 ;
  assign n25635 = n25625 ^ n25197 ;
  assign n25636 = ~n25624 & ~n25635 ;
  assign n25632 = n25346 ^ n24895 ;
  assign n25633 = n25632 ^ n24915 ;
  assign n25634 = n25633 ^ n25625 ;
  assign n25637 = n25636 ^ n25634 ;
  assign n25638 = n25637 ^ n25348 ;
  assign n25631 = n24749 ^ x344 ;
  assign n25639 = n25638 ^ n25631 ;
  assign n25628 = n25627 ^ n25619 ;
  assign n25629 = n25627 ^ n24749 ;
  assign n25630 = ~n25628 & ~n25629 ;
  assign n25640 = n25639 ^ n25630 ;
  assign n25885 = n25884 ^ n25640 ;
  assign n25995 = n25994 ^ n25885 ;
  assign n26003 = n25995 ^ n25014 ;
  assign n26004 = n26003 ^ n24456 ;
  assign n26005 = n25992 ^ n25002 ;
  assign n26006 = n26005 ^ n24387 ;
  assign n26007 = n25989 ^ n24990 ;
  assign n26008 = n26007 ^ n24366 ;
  assign n26009 = n25986 ^ n24978 ;
  assign n26010 = n26009 ^ n24345 ;
  assign n26011 = n25983 ^ n24955 ;
  assign n26012 = n26011 ^ n24320 ;
  assign n26014 = n25980 ^ n24952 ;
  assign n26087 = n25974 ^ n24901 ;
  assign n26015 = n25969 ^ n24885 ;
  assign n26016 = n26015 ^ n24086 ;
  assign n26017 = n25966 ^ n24864 ;
  assign n26018 = n26017 ^ n24166 ;
  assign n26019 = n25963 ^ n24843 ;
  assign n26020 = n26019 ^ n24160 ;
  assign n26075 = n26074 ^ n26072 ;
  assign n26076 = ~n26073 & ~n26075 ;
  assign n26077 = n26076 ^ n24154 ;
  assign n26078 = n26077 ^ n26019 ;
  assign n26079 = n26020 & ~n26078 ;
  assign n26080 = n26079 ^ n24160 ;
  assign n26081 = n26080 ^ n26017 ;
  assign n26082 = n26018 & ~n26081 ;
  assign n26083 = n26082 ^ n24166 ;
  assign n26084 = n26083 ^ n26015 ;
  assign n26085 = ~n26016 & n26084 ;
  assign n26086 = n26085 ^ n24086 ;
  assign n26088 = n26087 ^ n26086 ;
  assign n26089 = n25977 ^ n24923 ;
  assign n26090 = n26089 ^ n24181 ;
  assign n26091 = n26090 ^ n26086 ;
  assign n26092 = n26091 ^ n26089 ;
  assign n26093 = ~n26088 & ~n26092 ;
  assign n26094 = n26093 ^ n26090 ;
  assign n26097 = n25365 ^ n24285 ;
  assign n26098 = n26097 ^ n25980 ;
  assign n26095 = n25980 ^ n25365 ;
  assign n26096 = n26095 ^ n26089 ;
  assign n26099 = n26098 ^ n26096 ;
  assign n26100 = ~n26094 & n26099 ;
  assign n26101 = n26100 ^ n26098 ;
  assign n26102 = ~n26014 & n26101 ;
  assign n26013 = n26011 ^ n24300 ;
  assign n26103 = n26102 ^ n26013 ;
  assign n26104 = ~n26012 & n26103 ;
  assign n26105 = n26104 ^ n24320 ;
  assign n26106 = n26105 ^ n26009 ;
  assign n26107 = ~n26010 & ~n26106 ;
  assign n26108 = n26107 ^ n24345 ;
  assign n26109 = n26108 ^ n26007 ;
  assign n26110 = n26008 & ~n26109 ;
  assign n26111 = n26110 ^ n24366 ;
  assign n26112 = n26111 ^ n26005 ;
  assign n26113 = ~n26006 & ~n26112 ;
  assign n26114 = n26113 ^ n24387 ;
  assign n26115 = n26114 ^ n26003 ;
  assign n26116 = ~n26004 & ~n26115 ;
  assign n26117 = n26116 ^ n24456 ;
  assign n26135 = n26117 ^ n24488 ;
  assign n25998 = n25539 ^ n25528 ;
  assign n25996 = n25994 ^ n25528 ;
  assign n25997 = ~n25995 & ~n25996 ;
  assign n25999 = n25998 ^ n25997 ;
  assign n24939 = n24938 ^ x327 ;
  assign n26000 = n25999 ^ n24939 ;
  assign n26001 = n26000 ^ n25539 ;
  assign n26002 = n26001 ^ n25025 ;
  assign n26136 = n26135 ^ n26002 ;
  assign n26137 = n26136 ^ x432 ;
  assign n26234 = n26094 ^ n24285 ;
  assign n26138 = n26086 ^ n24181 ;
  assign n26139 = n26138 ^ n26087 ;
  assign n26140 = n26139 ^ x424 ;
  assign n26206 = n26077 ^ n24160 ;
  assign n26207 = n26206 ^ n26019 ;
  assign n26209 = n26207 ^ x428 ;
  assign n26208 = n26207 ^ n26200 ;
  assign n26210 = n26209 ^ n26208 ;
  assign n26211 = ~n26205 & n26210 ;
  assign n26212 = n26211 ^ n26209 ;
  assign n26213 = n26080 ^ n24166 ;
  assign n26214 = n26213 ^ n26017 ;
  assign n26216 = n26214 ^ x427 ;
  assign n26215 = n26214 ^ n26207 ;
  assign n26217 = n26216 ^ n26215 ;
  assign n26218 = ~n26212 & n26217 ;
  assign n26219 = n26218 ^ n26216 ;
  assign n26220 = n26083 ^ n24086 ;
  assign n26221 = n26220 ^ n26015 ;
  assign n26223 = n26221 ^ x426 ;
  assign n26222 = n26221 ^ n26214 ;
  assign n26224 = n26223 ^ n26222 ;
  assign n26225 = ~n26219 & n26224 ;
  assign n26226 = n26225 ^ n26223 ;
  assign n26228 = n26139 ^ x425 ;
  assign n26227 = n26221 ^ n26139 ;
  assign n26229 = n26228 ^ n26227 ;
  assign n26230 = n26226 & ~n26229 ;
  assign n26231 = n26230 ^ n26228 ;
  assign n26232 = ~n26140 & n26231 ;
  assign n26233 = n26232 ^ x424 ;
  assign n26235 = n26234 ^ n26233 ;
  assign n26236 = n26101 ^ n24300 ;
  assign n26237 = n26236 ^ x439 ;
  assign n26238 = n26237 ^ n26233 ;
  assign n26239 = n26238 ^ n26236 ;
  assign n26240 = n26235 & n26239 ;
  assign n26241 = n26240 ^ n26237 ;
  assign n26242 = n26103 ^ n24320 ;
  assign n26244 = n26242 ^ x438 ;
  assign n26243 = n26242 ^ n26236 ;
  assign n26245 = n26244 ^ n26243 ;
  assign n26246 = ~n26241 & n26245 ;
  assign n26247 = n26246 ^ n26244 ;
  assign n26248 = n26105 ^ n24345 ;
  assign n26249 = n26248 ^ n26009 ;
  assign n26251 = n26249 ^ x437 ;
  assign n26250 = n26249 ^ n26242 ;
  assign n26252 = n26251 ^ n26250 ;
  assign n26253 = ~n26247 & n26252 ;
  assign n26254 = n26253 ^ n26251 ;
  assign n26255 = n26108 ^ n24366 ;
  assign n26256 = n26255 ^ n26007 ;
  assign n26258 = n26256 ^ x436 ;
  assign n26257 = n26256 ^ n26249 ;
  assign n26259 = n26258 ^ n26257 ;
  assign n26260 = ~n26254 & n26259 ;
  assign n26261 = n26260 ^ n26258 ;
  assign n26262 = n26111 ^ n24387 ;
  assign n26263 = n26262 ^ n26005 ;
  assign n26265 = n26263 ^ x435 ;
  assign n26264 = n26263 ^ n26256 ;
  assign n26266 = n26265 ^ n26264 ;
  assign n26267 = ~n26261 & n26266 ;
  assign n26268 = n26267 ^ n26265 ;
  assign n26269 = n26114 ^ n24456 ;
  assign n26270 = n26269 ^ n26003 ;
  assign n26272 = n26270 ^ x434 ;
  assign n26271 = n26270 ^ n26263 ;
  assign n26273 = n26272 ^ n26271 ;
  assign n26274 = n26268 & ~n26273 ;
  assign n26275 = n26274 ^ n26272 ;
  assign n26277 = n26136 ^ x433 ;
  assign n26276 = n26270 ^ n26136 ;
  assign n26278 = n26277 ^ n26276 ;
  assign n26279 = ~n26275 & n26278 ;
  assign n26280 = n26279 ^ n26277 ;
  assign n26281 = n26137 & ~n26280 ;
  assign n26282 = n26281 ^ x432 ;
  assign n26118 = n26117 ^ n26002 ;
  assign n26124 = n25650 ^ x326 ;
  assign n26125 = n26124 ^ n25649 ;
  assign n26119 = n25548 ^ n25539 ;
  assign n26120 = n26119 ^ n25548 ;
  assign n26121 = n26120 ^ n24939 ;
  assign n26122 = ~n25999 & ~n26121 ;
  assign n26123 = n26122 ^ n26119 ;
  assign n26126 = n26125 ^ n26123 ;
  assign n26127 = n26126 ^ n25548 ;
  assign n26128 = n26127 ^ n25034 ;
  assign n26129 = n26128 ^ n24488 ;
  assign n26130 = n26129 ^ n26002 ;
  assign n26131 = n26130 ^ n26128 ;
  assign n26132 = ~n26118 & n26131 ;
  assign n26133 = n26132 ^ n26129 ;
  assign n26134 = n26133 ^ n24527 ;
  assign n26283 = n26282 ^ n26134 ;
  assign n26291 = n25560 ^ n24527 ;
  assign n26285 = n25658 ^ x325 ;
  assign n26287 = n26285 ^ n25548 ;
  assign n26286 = n26285 ^ n26125 ;
  assign n26288 = n26287 ^ n26286 ;
  assign n26289 = ~n26123 & n26288 ;
  assign n26290 = n26289 ^ n26287 ;
  assign n26292 = n26291 ^ n26290 ;
  assign n26284 = n26128 ^ n25560 ;
  assign n26293 = n26292 ^ n26284 ;
  assign n26294 = n26293 ^ n26290 ;
  assign n26295 = n26133 & ~n26294 ;
  assign n26296 = n26295 ^ n26292 ;
  assign n26297 = n26296 ^ n24562 ;
  assign n26298 = n26297 ^ x447 ;
  assign n26299 = n26298 ^ n26134 ;
  assign n26300 = n26299 ^ n26297 ;
  assign n26301 = n26283 & ~n26300 ;
  assign n26302 = n26301 ^ n26298 ;
  assign n26311 = n26290 ^ n25095 ;
  assign n26312 = n26296 & ~n26311 ;
  assign n26303 = n25665 ^ x324 ;
  assign n26305 = n26303 ^ n25561 ;
  assign n26304 = n26303 ^ n26285 ;
  assign n26306 = n26305 ^ n26304 ;
  assign n26307 = ~n26290 & n26306 ;
  assign n26308 = n26307 ^ n26305 ;
  assign n26309 = n26308 ^ n25114 ;
  assign n26310 = n26309 ^ n24562 ;
  assign n26313 = n26312 ^ n26310 ;
  assign n26314 = n26313 ^ n24595 ;
  assign n26316 = n26314 ^ x446 ;
  assign n26315 = n26314 ^ n26297 ;
  assign n26317 = n26316 ^ n26315 ;
  assign n26318 = n26302 & ~n26317 ;
  assign n26319 = n26318 ^ n26316 ;
  assign n26325 = n26303 ^ n25574 ;
  assign n26326 = n26308 & n26325 ;
  assign n26327 = n26326 ^ n25574 ;
  assign n26324 = n25833 ^ n25590 ;
  assign n26328 = n26327 ^ n26324 ;
  assign n26329 = n26328 ^ n25590 ;
  assign n26330 = n26329 ^ n25137 ;
  assign n26320 = n26309 ^ n24595 ;
  assign n26321 = ~n26313 & n26320 ;
  assign n26322 = n26321 ^ n24595 ;
  assign n26323 = n26322 ^ n24640 ;
  assign n26331 = n26330 ^ n26323 ;
  assign n26333 = n26331 ^ x445 ;
  assign n26332 = n26331 ^ n26314 ;
  assign n26334 = n26333 ^ n26332 ;
  assign n26335 = ~n26319 & n26334 ;
  assign n26336 = n26335 ^ n26333 ;
  assign n26348 = n25834 ^ n25833 ;
  assign n26342 = n26327 ^ n25590 ;
  assign n26345 = n26327 ^ n25833 ;
  assign n26346 = ~n26342 & n26345 ;
  assign n26343 = n25833 ^ n25602 ;
  assign n26347 = n26346 ^ n26343 ;
  assign n26349 = n26348 ^ n26347 ;
  assign n26350 = n26349 ^ n25602 ;
  assign n26351 = n26350 ^ n25157 ;
  assign n26337 = n26330 ^ n26322 ;
  assign n26338 = n26330 ^ n24640 ;
  assign n26339 = ~n26337 & ~n26338 ;
  assign n26340 = n26339 ^ n24640 ;
  assign n26341 = n26340 ^ n24681 ;
  assign n26352 = n26351 ^ n26341 ;
  assign n26354 = n26352 ^ x444 ;
  assign n26353 = n26352 ^ n26331 ;
  assign n26355 = n26354 ^ n26353 ;
  assign n26356 = n26336 & ~n26355 ;
  assign n26357 = n26356 ^ n26354 ;
  assign n26429 = n25836 ^ n25835 ;
  assign n26425 = n25614 ^ n25602 ;
  assign n26424 = n26348 ^ n25614 ;
  assign n26426 = n26425 ^ n26424 ;
  assign n26427 = ~n26347 & n26426 ;
  assign n26428 = n26427 ^ n26425 ;
  assign n26430 = n26429 ^ n26428 ;
  assign n26431 = n26430 ^ n25614 ;
  assign n26432 = n26431 ^ n25177 ;
  assign n26419 = n26351 ^ n26340 ;
  assign n26420 = n26351 ^ n24681 ;
  assign n26421 = ~n26419 & ~n26420 ;
  assign n26422 = n26421 ^ n24681 ;
  assign n26423 = n26422 ^ n24719 ;
  assign n26433 = n26432 ^ n26423 ;
  assign n26435 = n26433 ^ x443 ;
  assign n26434 = n26433 ^ n26352 ;
  assign n26436 = n26435 ^ n26434 ;
  assign n26437 = ~n26357 & n26436 ;
  assign n26438 = n26437 ^ n26435 ;
  assign n26439 = n26438 ^ x442 ;
  assign n26358 = n26357 ^ x443 ;
  assign n26380 = ~n26359 & n26379 ;
  assign n26381 = n26212 ^ x427 ;
  assign n26382 = n26380 & ~n26381 ;
  assign n26383 = n26219 ^ x426 ;
  assign n26384 = n26382 & ~n26383 ;
  assign n26385 = n26226 ^ x425 ;
  assign n26386 = n26384 & n26385 ;
  assign n26387 = n26231 ^ x424 ;
  assign n26388 = ~n26386 & ~n26387 ;
  assign n26389 = n26233 ^ x439 ;
  assign n26390 = n26389 ^ n26234 ;
  assign n26391 = ~n26388 & n26390 ;
  assign n26392 = n26241 ^ x438 ;
  assign n26393 = n26391 & ~n26392 ;
  assign n26394 = n26247 ^ x437 ;
  assign n26395 = ~n26393 & n26394 ;
  assign n26396 = n26254 ^ x436 ;
  assign n26397 = ~n26395 & ~n26396 ;
  assign n26398 = n26261 ^ x435 ;
  assign n26399 = n26397 & ~n26398 ;
  assign n26400 = n26268 ^ x434 ;
  assign n26401 = ~n26399 & ~n26400 ;
  assign n26402 = n26275 ^ x433 ;
  assign n26403 = n26401 & n26402 ;
  assign n26404 = n26280 ^ x432 ;
  assign n26405 = ~n26403 & ~n26404 ;
  assign n26406 = n26282 ^ x447 ;
  assign n26407 = n26406 ^ n26134 ;
  assign n26408 = ~n26405 & ~n26407 ;
  assign n26409 = n26302 ^ x446 ;
  assign n26410 = n26408 & ~n26409 ;
  assign n26411 = n26319 ^ x445 ;
  assign n26412 = n26410 & n26411 ;
  assign n26413 = n26336 ^ x444 ;
  assign n26414 = ~n26412 & n26413 ;
  assign n26440 = n26358 & ~n26414 ;
  assign n26478 = ~n26439 & ~n26440 ;
  assign n26464 = n25838 ^ n25837 ;
  assign n26466 = n26464 ^ n25614 ;
  assign n26465 = n26464 ^ n26429 ;
  assign n26467 = n26466 ^ n26465 ;
  assign n26468 = ~n26428 & ~n26467 ;
  assign n26469 = n26468 ^ n26466 ;
  assign n26470 = n26469 ^ n25197 ;
  assign n26459 = n26432 ^ n26422 ;
  assign n26460 = n26432 ^ n24719 ;
  assign n26461 = n26459 & n26460 ;
  assign n26462 = n26461 ^ n24719 ;
  assign n26463 = n26462 ^ n24756 ;
  assign n26471 = n26470 ^ n26463 ;
  assign n26473 = n26471 ^ x442 ;
  assign n26472 = n26471 ^ n26433 ;
  assign n26474 = n26473 ^ n26472 ;
  assign n26475 = ~n26438 & n26474 ;
  assign n26476 = n26475 ^ n26473 ;
  assign n26477 = n26476 ^ x441 ;
  assign n26479 = n26478 ^ n26477 ;
  assign n26498 = n26497 ^ n26479 ;
  assign n26456 = n25930 ^ n25407 ;
  assign n26457 = n26456 ^ n25921 ;
  assign n26444 = n25927 ^ n25926 ;
  assign n26415 = n26414 ^ n26358 ;
  assign n26442 = n25924 ^ n25923 ;
  assign n26443 = ~n26415 & n26442 ;
  assign n26445 = n26444 ^ n26443 ;
  assign n26441 = n26440 ^ n26439 ;
  assign n26453 = n26443 ^ n26441 ;
  assign n26454 = ~n26445 & n26453 ;
  assign n26455 = n26454 ^ n26444 ;
  assign n26458 = n26457 ^ n26455 ;
  assign n26494 = n26479 ^ n26457 ;
  assign n26495 = n26458 & ~n26494 ;
  assign n26499 = n26498 ^ n26495 ;
  assign n26516 = n26478 ^ n26471 ;
  assign n26519 = ~n26476 & n26516 ;
  assign n26515 = n26476 ^ n26471 ;
  assign n26517 = n26516 ^ n26515 ;
  assign n26518 = ~x441 & ~n26517 ;
  assign n26520 = n26519 ^ n26518 ;
  assign n26507 = n26464 ^ n25626 ;
  assign n26508 = ~n26469 & ~n26507 ;
  assign n26504 = n25839 ^ n25637 ;
  assign n26505 = n26504 ^ n25840 ;
  assign n26506 = n26505 ^ n26464 ;
  assign n26509 = n26508 ^ n26506 ;
  assign n26510 = n26509 ^ n25637 ;
  assign n26511 = n26510 ^ n25346 ;
  assign n26512 = n26511 ^ n24795 ;
  assign n26503 = n24756 ^ x440 ;
  assign n26513 = n26512 ^ n26503 ;
  assign n26500 = n26470 ^ n26462 ;
  assign n26501 = n26470 ^ n24756 ;
  assign n26502 = n26500 & ~n26501 ;
  assign n26514 = n26513 ^ n26502 ;
  assign n26521 = n26520 ^ n26514 ;
  assign n26536 = n26521 ^ n26497 ;
  assign n26537 = n26499 & ~n26536 ;
  assign n26540 = n26539 ^ n26537 ;
  assign n26541 = n26144 ^ x423 ;
  assign n26556 = n26541 ^ n26538 ;
  assign n26557 = ~n26540 & ~n26556 ;
  assign n26558 = n26557 ^ n26541 ;
  assign n26576 = n26560 ^ n26558 ;
  assign n26577 = n25944 ^ n25429 ;
  assign n26578 = n26577 ^ n25915 ;
  assign n26579 = n26578 ^ n26361 ;
  assign n26580 = n26579 ^ n26578 ;
  assign n26581 = n26580 ^ n26558 ;
  assign n26582 = ~n26576 & n26581 ;
  assign n26583 = n26582 ^ n26579 ;
  assign n26584 = n25947 ^ n25435 ;
  assign n26585 = n26584 ^ n25913 ;
  assign n26588 = n26585 ^ n26578 ;
  assign n26586 = n26362 ^ n26361 ;
  assign n26587 = n26586 ^ n26585 ;
  assign n26589 = n26588 ^ n26587 ;
  assign n26590 = ~n26583 & n26589 ;
  assign n26591 = n26590 ^ n26588 ;
  assign n26592 = n25950 ^ n25441 ;
  assign n26593 = n26592 ^ n25911 ;
  assign n26596 = n26593 ^ n26585 ;
  assign n26594 = n26364 ^ n26363 ;
  assign n26595 = n26594 ^ n26593 ;
  assign n26597 = n26596 ^ n26595 ;
  assign n26598 = ~n26591 & n26597 ;
  assign n26599 = n26598 ^ n26596 ;
  assign n26600 = n25953 ^ n25447 ;
  assign n26601 = n26600 ^ n25909 ;
  assign n26604 = n26601 ^ n26593 ;
  assign n26602 = n26366 ^ n26365 ;
  assign n26603 = n26602 ^ n26601 ;
  assign n26605 = n26604 ^ n26603 ;
  assign n26606 = ~n26599 & n26605 ;
  assign n26607 = n26606 ^ n26604 ;
  assign n26608 = n25956 ^ n25453 ;
  assign n26609 = n26608 ^ n25907 ;
  assign n26612 = n26609 ^ n26601 ;
  assign n26610 = n26368 ^ n26367 ;
  assign n26611 = n26610 ^ n26609 ;
  assign n26613 = n26612 ^ n26611 ;
  assign n26614 = ~n26607 & n26613 ;
  assign n26615 = n26614 ^ n26612 ;
  assign n26616 = n25959 ^ n25459 ;
  assign n26617 = n26616 ^ n25905 ;
  assign n26620 = n26617 ^ n26609 ;
  assign n26618 = n26370 ^ n26369 ;
  assign n26619 = n26618 ^ n26617 ;
  assign n26621 = n26620 ^ n26619 ;
  assign n26622 = n26615 & n26621 ;
  assign n26623 = n26622 ^ n26620 ;
  assign n26624 = n25962 ^ n25466 ;
  assign n26625 = n26624 ^ n25903 ;
  assign n26628 = n26625 ^ n26617 ;
  assign n26626 = n26372 ^ n26371 ;
  assign n26627 = n26626 ^ n26625 ;
  assign n26629 = n26628 ^ n26627 ;
  assign n26630 = n26623 & ~n26629 ;
  assign n26631 = n26630 ^ n26628 ;
  assign n26632 = n25965 ^ n25472 ;
  assign n26633 = n26632 ^ n25901 ;
  assign n26636 = n26633 ^ n26625 ;
  assign n26634 = n26374 ^ n26373 ;
  assign n26635 = n26634 ^ n26633 ;
  assign n26637 = n26636 ^ n26635 ;
  assign n26638 = ~n26631 & n26637 ;
  assign n26639 = n26638 ^ n26636 ;
  assign n26640 = n25968 ^ n25393 ;
  assign n26641 = n26640 ^ n25899 ;
  assign n26644 = n26641 ^ n26633 ;
  assign n26642 = n26376 ^ n26375 ;
  assign n26643 = n26642 ^ n26641 ;
  assign n26645 = n26644 ^ n26643 ;
  assign n26646 = ~n26639 & n26645 ;
  assign n26647 = n26646 ^ n26644 ;
  assign n26648 = n25973 ^ n25972 ;
  assign n26651 = n26648 ^ n26641 ;
  assign n26649 = n26378 ^ n26377 ;
  assign n26650 = n26649 ^ n26648 ;
  assign n26652 = n26651 ^ n26650 ;
  assign n26653 = ~n26647 & n26652 ;
  assign n26654 = n26653 ^ n26651 ;
  assign n26656 = n26655 ^ n26654 ;
  assign n26416 = n26415 ^ n24937 ;
  assign n26448 = n25244 & n26416 ;
  assign n26446 = n26445 ^ n26441 ;
  assign n26447 = n26446 ^ n25928 ;
  assign n26449 = n26448 ^ n26447 ;
  assign n26450 = n26449 ^ n25246 ;
  assign n26417 = x7 & ~n26416 ;
  assign n26452 = n26450 ^ n26417 ;
  assign n26482 = n26448 ^ n25246 ;
  assign n26483 = ~n26449 & ~n26482 ;
  assign n26484 = n26483 ^ n25246 ;
  assign n26485 = n26484 ^ n25248 ;
  assign n26480 = n26479 ^ n26458 ;
  assign n26481 = n26480 ^ n25931 ;
  assign n26486 = n26485 ^ n26481 ;
  assign n26487 = n26486 ^ x6 ;
  assign n26488 = n26487 ^ n26450 ;
  assign n26489 = n26488 ^ n26486 ;
  assign n26490 = n26452 & ~n26489 ;
  assign n26491 = n26490 ^ n26487 ;
  assign n26524 = n26484 ^ n26481 ;
  assign n26525 = n26485 & n26524 ;
  assign n26526 = n26525 ^ n25248 ;
  assign n26527 = n26526 ^ n25256 ;
  assign n26522 = n26521 ^ n26499 ;
  assign n26523 = n26522 ^ n25934 ;
  assign n26528 = n26527 ^ n26523 ;
  assign n26530 = n26528 ^ x5 ;
  assign n26529 = n26528 ^ n26486 ;
  assign n26531 = n26530 ^ n26529 ;
  assign n26532 = ~n26491 & n26531 ;
  assign n26533 = n26532 ^ n26530 ;
  assign n26544 = n26526 ^ n26523 ;
  assign n26545 = ~n26527 & n26544 ;
  assign n26546 = n26545 ^ n25256 ;
  assign n26547 = n26546 ^ n25264 ;
  assign n26542 = n26541 ^ n26540 ;
  assign n26543 = n26542 ^ n25939 ;
  assign n26548 = n26547 ^ n26543 ;
  assign n26550 = n26548 ^ x4 ;
  assign n26549 = n26548 ^ n26528 ;
  assign n26551 = n26550 ^ n26549 ;
  assign n26552 = n26533 & ~n26551 ;
  assign n26553 = n26552 ^ n26550 ;
  assign n26554 = n26553 ^ x3 ;
  assign n26418 = n26417 ^ x6 ;
  assign n26451 = n26450 ^ n26418 ;
  assign n26492 = n26491 ^ x5 ;
  assign n26493 = ~n26451 & n26492 ;
  assign n26534 = n26533 ^ x4 ;
  assign n26535 = ~n26493 & n26534 ;
  assign n26575 = n26554 ^ n26535 ;
  assign n26657 = n26656 ^ n26575 ;
  assign n26811 = n26394 ^ n26393 ;
  assign n26668 = n26383 ^ n26382 ;
  assign n26660 = n26381 ^ n26380 ;
  assign n26658 = n25976 ^ n25483 ;
  assign n26659 = n26658 ^ n25897 ;
  assign n26661 = n26660 ^ n26659 ;
  assign n26662 = n26655 ^ n26648 ;
  assign n26663 = n26654 & ~n26662 ;
  assign n26664 = n26663 ^ n26648 ;
  assign n26665 = n26664 ^ n26660 ;
  assign n26666 = ~n26661 & ~n26665 ;
  assign n26667 = n26666 ^ n26664 ;
  assign n26669 = n26668 ^ n26667 ;
  assign n26672 = n25979 ^ n25490 ;
  assign n26673 = n26672 ^ n25895 ;
  assign n26676 = n26673 ^ n26667 ;
  assign n26677 = n26669 & ~n26676 ;
  assign n26670 = n25982 ^ n25389 ;
  assign n26671 = n26670 ^ n25893 ;
  assign n26674 = n26673 ^ n26671 ;
  assign n26678 = n26677 ^ n26674 ;
  assign n26763 = n25985 ^ n25386 ;
  assign n26764 = n26763 ^ n25891 ;
  assign n26766 = n26764 ^ n26671 ;
  assign n26679 = n26385 ^ n26384 ;
  assign n26765 = n26764 ^ n26679 ;
  assign n26767 = n26766 ^ n26765 ;
  assign n26768 = ~n26678 & n26767 ;
  assign n26769 = n26768 ^ n26766 ;
  assign n26777 = n25988 ^ n25383 ;
  assign n26778 = n26777 ^ n25889 ;
  assign n26780 = n26778 ^ n26764 ;
  assign n26770 = n26387 ^ n26386 ;
  assign n26779 = n26778 ^ n26770 ;
  assign n26781 = n26780 ^ n26779 ;
  assign n26782 = ~n26769 & n26781 ;
  assign n26783 = n26782 ^ n26780 ;
  assign n26791 = n25991 ^ n25515 ;
  assign n26792 = n26791 ^ n25887 ;
  assign n26794 = n26792 ^ n26778 ;
  assign n26784 = n26390 ^ n26388 ;
  assign n26793 = n26792 ^ n26784 ;
  assign n26795 = n26794 ^ n26793 ;
  assign n26796 = ~n26783 & ~n26795 ;
  assign n26797 = n26796 ^ n26794 ;
  assign n26805 = n25996 ^ n25885 ;
  assign n26807 = n26805 ^ n26792 ;
  assign n26798 = n26392 ^ n26391 ;
  assign n26806 = n26805 ^ n26798 ;
  assign n26808 = n26807 ^ n26806 ;
  assign n26809 = ~n26797 & n26808 ;
  assign n26810 = n26809 ^ n26807 ;
  assign n26812 = n26811 ^ n26810 ;
  assign n26813 = n26812 ^ n25995 ;
  assign n26799 = n26798 ^ n26797 ;
  assign n26800 = n26799 ^ n25992 ;
  assign n26785 = n26784 ^ n26783 ;
  assign n26786 = n26785 ^ n25989 ;
  assign n26771 = n26770 ^ n26769 ;
  assign n26772 = n26771 ^ n25986 ;
  assign n26680 = n26679 ^ n26678 ;
  assign n26681 = n26680 ^ n25983 ;
  assign n26682 = n26681 ^ n24955 ;
  assign n26684 = n26586 ^ n26583 ;
  assign n26685 = n26684 ^ n25945 ;
  assign n26686 = n26685 ^ n25279 ;
  assign n26564 = n26546 ^ n26543 ;
  assign n26565 = n26547 & n26564 ;
  assign n26566 = n26565 ^ n25264 ;
  assign n26567 = n26566 ^ n25271 ;
  assign n26561 = n26560 ^ n26361 ;
  assign n26562 = n26561 ^ n26558 ;
  assign n26563 = n26562 ^ n25942 ;
  assign n26687 = n26566 ^ n26563 ;
  assign n26688 = n26567 & n26687 ;
  assign n26689 = n26688 ^ n25271 ;
  assign n26690 = n26689 ^ n26685 ;
  assign n26691 = n26686 & ~n26690 ;
  assign n26692 = n26691 ^ n25279 ;
  assign n26693 = n26692 ^ n25287 ;
  assign n26694 = n26594 ^ n26591 ;
  assign n26695 = n26694 ^ n25948 ;
  assign n26696 = n26695 ^ n26692 ;
  assign n26697 = n26693 & n26696 ;
  assign n26698 = n26697 ^ n25287 ;
  assign n26699 = n26698 ^ n25295 ;
  assign n26700 = n26602 ^ n26599 ;
  assign n26701 = n26700 ^ n25951 ;
  assign n26702 = n26701 ^ n26698 ;
  assign n26703 = ~n26699 & n26702 ;
  assign n26704 = n26703 ^ n25295 ;
  assign n26705 = n26704 ^ n25302 ;
  assign n26706 = n26610 ^ n26607 ;
  assign n26707 = n26706 ^ n25954 ;
  assign n26708 = n26707 ^ n26704 ;
  assign n26709 = n26705 & ~n26708 ;
  assign n26710 = n26709 ^ n25302 ;
  assign n26711 = n26710 ^ n25310 ;
  assign n26712 = n26618 ^ n26615 ;
  assign n26713 = n26712 ^ n25957 ;
  assign n26714 = n26713 ^ n26710 ;
  assign n26715 = ~n26711 & n26714 ;
  assign n26716 = n26715 ^ n25310 ;
  assign n26717 = n26716 ^ n25242 ;
  assign n26718 = n26626 ^ n26623 ;
  assign n26719 = n26718 ^ n25960 ;
  assign n26720 = n26719 ^ n26716 ;
  assign n26721 = ~n26717 & n26720 ;
  assign n26722 = n26721 ^ n25242 ;
  assign n26723 = n26722 ^ n24843 ;
  assign n26724 = n26634 ^ n26631 ;
  assign n26725 = n26724 ^ n25963 ;
  assign n26726 = n26725 ^ n26722 ;
  assign n26727 = ~n26723 & n26726 ;
  assign n26728 = n26727 ^ n24843 ;
  assign n26729 = n26728 ^ n24864 ;
  assign n26730 = n26642 ^ n26639 ;
  assign n26731 = n26730 ^ n25966 ;
  assign n26732 = n26731 ^ n26728 ;
  assign n26733 = ~n26729 & ~n26732 ;
  assign n26734 = n26733 ^ n24864 ;
  assign n26735 = n26734 ^ n24885 ;
  assign n26736 = n26649 ^ n26647 ;
  assign n26737 = n26736 ^ n25969 ;
  assign n26738 = n26737 ^ n26734 ;
  assign n26739 = n26735 & n26738 ;
  assign n26740 = n26739 ^ n24885 ;
  assign n26683 = n26656 ^ n25974 ;
  assign n26741 = n26740 ^ n26683 ;
  assign n26742 = n26664 ^ n26661 ;
  assign n26743 = n26742 ^ n25977 ;
  assign n26744 = n26743 ^ n24901 ;
  assign n26745 = n26744 ^ n26683 ;
  assign n26746 = n26745 ^ n26743 ;
  assign n26747 = n26741 & n26746 ;
  assign n26748 = n26747 ^ n26744 ;
  assign n26749 = n26673 ^ n26669 ;
  assign n26750 = n26749 ^ n25980 ;
  assign n26752 = n26750 ^ n24923 ;
  assign n26751 = n26750 ^ n26743 ;
  assign n26753 = n26752 ^ n26751 ;
  assign n26754 = n26748 & n26753 ;
  assign n26755 = n26754 ^ n26752 ;
  assign n26757 = n26681 ^ n25365 ;
  assign n26756 = n26750 ^ n26681 ;
  assign n26758 = n26757 ^ n26756 ;
  assign n26759 = ~n26755 & ~n26758 ;
  assign n26760 = n26759 ^ n26757 ;
  assign n26761 = n26682 & ~n26760 ;
  assign n26762 = n26761 ^ n24955 ;
  assign n26773 = n26772 ^ n26762 ;
  assign n26774 = n26772 ^ n24978 ;
  assign n26775 = n26773 & n26774 ;
  assign n26776 = n26775 ^ n24978 ;
  assign n26787 = n26786 ^ n26776 ;
  assign n26788 = n26786 ^ n24990 ;
  assign n26789 = n26787 & ~n26788 ;
  assign n26790 = n26789 ^ n24990 ;
  assign n26801 = n26800 ^ n26790 ;
  assign n26802 = n26800 ^ n25002 ;
  assign n26803 = ~n26801 & ~n26802 ;
  assign n26804 = n26803 ^ n25002 ;
  assign n26814 = n26813 ^ n26804 ;
  assign n26815 = n26813 ^ n25014 ;
  assign n26816 = ~n26814 & ~n26815 ;
  assign n26817 = n26816 ^ n25014 ;
  assign n26839 = n26817 ^ n25025 ;
  assign n26820 = n26811 ^ n26805 ;
  assign n26821 = ~n26810 & n26820 ;
  assign n26819 = n26805 ^ n26000 ;
  assign n26822 = n26821 ^ n26819 ;
  assign n26818 = n26396 ^ n26395 ;
  assign n26823 = n26822 ^ n26818 ;
  assign n26824 = n26823 ^ n26001 ;
  assign n26840 = n26839 ^ n26824 ;
  assign n26841 = n26840 ^ x16 ;
  assign n26843 = n26740 ^ n24901 ;
  assign n26844 = n26843 ^ n26683 ;
  assign n26845 = n26844 ^ x8 ;
  assign n26569 = n26548 ^ x3 ;
  assign n26570 = n26553 & ~n26569 ;
  assign n26571 = n26570 ^ x3 ;
  assign n26568 = n26567 ^ n26563 ;
  assign n26572 = n26571 ^ n26568 ;
  assign n26848 = n26571 ^ x2 ;
  assign n26849 = n26572 & n26848 ;
  assign n26850 = n26849 ^ x2 ;
  assign n26846 = n26689 ^ n25279 ;
  assign n26847 = n26846 ^ n26685 ;
  assign n26851 = n26850 ^ n26847 ;
  assign n26852 = n26695 ^ n26693 ;
  assign n26853 = n26852 ^ x1 ;
  assign n26854 = n26853 ^ n26850 ;
  assign n26855 = n26854 ^ n26852 ;
  assign n26856 = ~n26851 & n26855 ;
  assign n26857 = n26856 ^ n26853 ;
  assign n26858 = n26701 ^ n26699 ;
  assign n26860 = n26858 ^ x0 ;
  assign n26859 = n26858 ^ n26852 ;
  assign n26861 = n26860 ^ n26859 ;
  assign n26862 = n26857 & ~n26861 ;
  assign n26863 = n26862 ^ n26860 ;
  assign n26864 = n26707 ^ n26705 ;
  assign n26866 = n26864 ^ x15 ;
  assign n26865 = n26864 ^ n26858 ;
  assign n26867 = n26866 ^ n26865 ;
  assign n26868 = ~n26863 & n26867 ;
  assign n26869 = n26868 ^ n26866 ;
  assign n26870 = n26713 ^ n26711 ;
  assign n26872 = n26870 ^ x14 ;
  assign n26871 = n26870 ^ n26864 ;
  assign n26873 = n26872 ^ n26871 ;
  assign n26874 = n26869 & ~n26873 ;
  assign n26875 = n26874 ^ n26872 ;
  assign n26876 = n26719 ^ n26717 ;
  assign n26878 = n26876 ^ x13 ;
  assign n26877 = n26876 ^ n26870 ;
  assign n26879 = n26878 ^ n26877 ;
  assign n26880 = n26875 & ~n26879 ;
  assign n26881 = n26880 ^ n26878 ;
  assign n26882 = n26725 ^ n26723 ;
  assign n26884 = n26882 ^ x12 ;
  assign n26883 = n26882 ^ n26876 ;
  assign n26885 = n26884 ^ n26883 ;
  assign n26886 = ~n26881 & n26885 ;
  assign n26887 = n26886 ^ n26884 ;
  assign n26888 = n26731 ^ n26729 ;
  assign n26890 = n26888 ^ x11 ;
  assign n26889 = n26888 ^ n26882 ;
  assign n26891 = n26890 ^ n26889 ;
  assign n26892 = n26887 & ~n26891 ;
  assign n26893 = n26892 ^ n26890 ;
  assign n26894 = n26737 ^ n26735 ;
  assign n26896 = n26894 ^ x10 ;
  assign n26895 = n26894 ^ n26888 ;
  assign n26897 = n26896 ^ n26895 ;
  assign n26898 = n26893 & ~n26897 ;
  assign n26899 = n26898 ^ n26896 ;
  assign n26901 = n26844 ^ x9 ;
  assign n26900 = n26894 ^ n26844 ;
  assign n26902 = n26901 ^ n26900 ;
  assign n26903 = ~n26899 & n26902 ;
  assign n26904 = n26903 ^ n26901 ;
  assign n26905 = ~n26845 & n26904 ;
  assign n26906 = n26905 ^ x8 ;
  assign n26842 = n26748 ^ n24923 ;
  assign n26907 = n26906 ^ n26842 ;
  assign n26908 = n26755 ^ n25365 ;
  assign n26909 = n26908 ^ x23 ;
  assign n26910 = n26909 ^ n26842 ;
  assign n26911 = n26910 ^ n26908 ;
  assign n26912 = ~n26907 & n26911 ;
  assign n26913 = n26912 ^ n26909 ;
  assign n26914 = n26760 ^ n24955 ;
  assign n26916 = n26914 ^ x22 ;
  assign n26915 = n26914 ^ n26908 ;
  assign n26917 = n26916 ^ n26915 ;
  assign n26918 = ~n26913 & n26917 ;
  assign n26919 = n26918 ^ n26916 ;
  assign n26920 = n26762 ^ n24978 ;
  assign n26921 = n26920 ^ n26772 ;
  assign n26923 = n26921 ^ x21 ;
  assign n26922 = n26921 ^ n26914 ;
  assign n26924 = n26923 ^ n26922 ;
  assign n26925 = ~n26919 & n26924 ;
  assign n26926 = n26925 ^ n26923 ;
  assign n26927 = n26776 ^ n24990 ;
  assign n26928 = n26927 ^ n26786 ;
  assign n26930 = n26928 ^ x20 ;
  assign n26929 = n26928 ^ n26921 ;
  assign n26931 = n26930 ^ n26929 ;
  assign n26932 = ~n26926 & n26931 ;
  assign n26933 = n26932 ^ n26930 ;
  assign n26934 = n26790 ^ n25002 ;
  assign n26935 = n26934 ^ n26800 ;
  assign n26937 = n26935 ^ x19 ;
  assign n26936 = n26935 ^ n26928 ;
  assign n26938 = n26937 ^ n26936 ;
  assign n26939 = ~n26933 & n26938 ;
  assign n26940 = n26939 ^ n26937 ;
  assign n26941 = n26804 ^ n25014 ;
  assign n26942 = n26941 ^ n26813 ;
  assign n26944 = n26942 ^ x18 ;
  assign n26943 = n26942 ^ n26935 ;
  assign n26945 = n26944 ^ n26943 ;
  assign n26946 = ~n26940 & n26945 ;
  assign n26947 = n26946 ^ n26944 ;
  assign n26949 = n26840 ^ x17 ;
  assign n26948 = n26942 ^ n26840 ;
  assign n26950 = n26949 ^ n26948 ;
  assign n26951 = n26947 & ~n26950 ;
  assign n26952 = n26951 ^ n26949 ;
  assign n26953 = ~n26841 & n26952 ;
  assign n26954 = n26953 ^ x16 ;
  assign n26825 = n26824 ^ n26817 ;
  assign n26828 = n26818 ^ n26000 ;
  assign n26829 = ~n26822 & ~n26828 ;
  assign n26830 = n26829 ^ n26000 ;
  assign n26826 = n26398 ^ n26397 ;
  assign n26827 = n26826 ^ n26126 ;
  assign n26831 = n26830 ^ n26827 ;
  assign n26832 = n26831 ^ n26127 ;
  assign n26833 = n26832 ^ n25025 ;
  assign n26834 = n26833 ^ n26832 ;
  assign n26835 = n26834 ^ n26817 ;
  assign n26836 = n26825 & ~n26835 ;
  assign n26837 = n26836 ^ n26833 ;
  assign n26838 = n26837 ^ n25034 ;
  assign n26955 = n26954 ^ n26838 ;
  assign n26962 = n26290 ^ n25561 ;
  assign n26960 = n26400 ^ n26399 ;
  assign n26956 = n26830 ^ n26826 ;
  assign n26957 = n26830 ^ n26126 ;
  assign n26958 = ~n26956 & n26957 ;
  assign n26959 = n26958 ^ n26126 ;
  assign n26961 = n26960 ^ n26959 ;
  assign n26963 = n26962 ^ n26961 ;
  assign n26964 = n26963 ^ n26290 ;
  assign n26966 = n26964 ^ n25034 ;
  assign n26965 = n26964 ^ n26832 ;
  assign n26967 = n26966 ^ n26965 ;
  assign n26968 = n26837 & ~n26967 ;
  assign n26969 = n26968 ^ n26966 ;
  assign n26970 = n26969 ^ n25560 ;
  assign n26971 = n26970 ^ x31 ;
  assign n26972 = n26971 ^ n26838 ;
  assign n26973 = n26972 ^ n26970 ;
  assign n26974 = n26955 & ~n26973 ;
  assign n26975 = n26974 ^ n26971 ;
  assign n26982 = n26402 ^ n26401 ;
  assign n26976 = n26308 ^ n25574 ;
  assign n26977 = n26976 ^ n26962 ;
  assign n26978 = n26977 ^ n26960 ;
  assign n26979 = n26978 ^ n26976 ;
  assign n26980 = ~n26961 & ~n26979 ;
  assign n26981 = n26980 ^ n26977 ;
  assign n26983 = n26982 ^ n26981 ;
  assign n26984 = n26983 ^ n26308 ;
  assign n26986 = n26984 ^ n25560 ;
  assign n26985 = n26984 ^ n26964 ;
  assign n26987 = n26986 ^ n26985 ;
  assign n26988 = n26969 & n26987 ;
  assign n26989 = n26988 ^ n26986 ;
  assign n26990 = n26989 ^ n25114 ;
  assign n26992 = n26990 ^ x30 ;
  assign n26991 = n26990 ^ n26970 ;
  assign n26993 = n26992 ^ n26991 ;
  assign n26994 = ~n26975 & n26993 ;
  assign n26995 = n26994 ^ n26992 ;
  assign n27002 = n26982 ^ n26976 ;
  assign n27003 = n26981 & ~n27002 ;
  assign n27001 = n26976 ^ n26328 ;
  assign n27004 = n27003 ^ n27001 ;
  assign n27000 = n26404 ^ n26403 ;
  assign n27005 = n27004 ^ n27000 ;
  assign n27006 = n27005 ^ n26329 ;
  assign n26996 = n26984 ^ n25114 ;
  assign n26997 = ~n26989 & n26996 ;
  assign n26998 = n26997 ^ n25114 ;
  assign n26999 = n26998 ^ n25137 ;
  assign n27007 = n27006 ^ n26999 ;
  assign n27009 = n27007 ^ x29 ;
  assign n27008 = n27007 ^ n26990 ;
  assign n27010 = n27009 ^ n27008 ;
  assign n27011 = n26995 & ~n27010 ;
  assign n27012 = n27011 ^ n27009 ;
  assign n27023 = n26407 ^ n26405 ;
  assign n27018 = n26349 ^ n26328 ;
  assign n27019 = n27018 ^ n26349 ;
  assign n27020 = n27019 ^ n27000 ;
  assign n27021 = ~n27004 & ~n27020 ;
  assign n27022 = n27021 ^ n27018 ;
  assign n27024 = n27023 ^ n27022 ;
  assign n27025 = n27024 ^ n26350 ;
  assign n27013 = n27006 ^ n26998 ;
  assign n27014 = n27006 ^ n25137 ;
  assign n27015 = n27013 & n27014 ;
  assign n27016 = n27015 ^ n25137 ;
  assign n27017 = n27016 ^ n25157 ;
  assign n27026 = n27025 ^ n27017 ;
  assign n27028 = n27026 ^ x28 ;
  assign n27027 = n27026 ^ n27007 ;
  assign n27029 = n27028 ^ n27027 ;
  assign n27030 = n27012 & ~n27029 ;
  assign n27031 = n27030 ^ n27028 ;
  assign n27042 = n26409 ^ n26408 ;
  assign n27038 = n26430 ^ n26349 ;
  assign n27037 = n27023 ^ n26430 ;
  assign n27039 = n27038 ^ n27037 ;
  assign n27040 = n27022 & n27039 ;
  assign n27041 = n27040 ^ n27038 ;
  assign n27043 = n27042 ^ n27041 ;
  assign n27044 = n27043 ^ n26431 ;
  assign n27032 = n27025 ^ n27016 ;
  assign n27033 = n27025 ^ n25157 ;
  assign n27034 = n27032 & ~n27033 ;
  assign n27035 = n27034 ^ n25157 ;
  assign n27036 = n27035 ^ n25177 ;
  assign n27045 = n27044 ^ n27036 ;
  assign n27047 = n27045 ^ x27 ;
  assign n27046 = n27045 ^ n27026 ;
  assign n27048 = n27047 ^ n27046 ;
  assign n27049 = n27031 & ~n27048 ;
  assign n27050 = n27049 ^ n27047 ;
  assign n27113 = n26411 ^ n26410 ;
  assign n27107 = n26469 ^ n25626 ;
  assign n27109 = n27107 ^ n26430 ;
  assign n27108 = n27107 ^ n27042 ;
  assign n27110 = n27109 ^ n27108 ;
  assign n27111 = n27041 & ~n27110 ;
  assign n27112 = n27111 ^ n27109 ;
  assign n27114 = n27113 ^ n27112 ;
  assign n27115 = n27114 ^ n26469 ;
  assign n27102 = n27044 ^ n27035 ;
  assign n27103 = n27044 ^ n25177 ;
  assign n27104 = n27102 & n27103 ;
  assign n27105 = n27104 ^ n25177 ;
  assign n27106 = n27105 ^ n25197 ;
  assign n27116 = n27115 ^ n27106 ;
  assign n27118 = n27116 ^ x26 ;
  assign n27117 = n27116 ^ n27045 ;
  assign n27119 = n27118 ^ n27117 ;
  assign n27120 = ~n27050 & n27119 ;
  assign n27121 = n27120 ^ n27118 ;
  assign n27051 = n27050 ^ x26 ;
  assign n27052 = n27031 ^ x27 ;
  assign n27053 = n26995 ^ x29 ;
  assign n27054 = n26975 ^ x30 ;
  assign n27055 = n26954 ^ x31 ;
  assign n27056 = n27055 ^ n26838 ;
  assign n27057 = n26952 ^ x16 ;
  assign n27058 = n26947 ^ x17 ;
  assign n27059 = n26940 ^ x18 ;
  assign n26555 = n26535 & n26554 ;
  assign n26573 = n26572 ^ x2 ;
  assign n27060 = n26555 & n26573 ;
  assign n27061 = n26851 ^ x1 ;
  assign n27062 = n27060 & ~n27061 ;
  assign n27063 = n26857 ^ x0 ;
  assign n27064 = n27062 & n27063 ;
  assign n27065 = n26863 ^ x15 ;
  assign n27066 = n27064 & ~n27065 ;
  assign n27067 = n26869 ^ x14 ;
  assign n27068 = n27066 & n27067 ;
  assign n27069 = n26875 ^ x13 ;
  assign n27070 = n27068 & n27069 ;
  assign n27071 = n26881 ^ x12 ;
  assign n27072 = ~n27070 & n27071 ;
  assign n27073 = n26887 ^ x11 ;
  assign n27074 = n27072 & ~n27073 ;
  assign n27075 = n26893 ^ x10 ;
  assign n27076 = ~n27074 & n27075 ;
  assign n27077 = n26899 ^ x9 ;
  assign n27078 = ~n27076 & n27077 ;
  assign n27079 = n26904 ^ x8 ;
  assign n27080 = n27078 & ~n27079 ;
  assign n27081 = n26906 ^ x23 ;
  assign n27082 = n27081 ^ n26842 ;
  assign n27083 = ~n27080 & ~n27082 ;
  assign n27084 = n26913 ^ x22 ;
  assign n27085 = ~n27083 & n27084 ;
  assign n27086 = n26919 ^ x21 ;
  assign n27087 = n27085 & n27086 ;
  assign n27088 = n26926 ^ x20 ;
  assign n27089 = n27087 & n27088 ;
  assign n27090 = n26933 ^ x19 ;
  assign n27091 = n27089 & n27090 ;
  assign n27092 = ~n27059 & ~n27091 ;
  assign n27093 = ~n27058 & ~n27092 ;
  assign n27094 = n27057 & ~n27093 ;
  assign n27095 = ~n27056 & ~n27094 ;
  assign n27096 = ~n27054 & ~n27095 ;
  assign n27097 = ~n27053 & ~n27096 ;
  assign n27098 = n27012 ^ x28 ;
  assign n27099 = ~n27097 & n27098 ;
  assign n27100 = ~n27052 & ~n27099 ;
  assign n27101 = ~n27051 & ~n27100 ;
  assign n27185 = n27116 ^ n27101 ;
  assign n27188 = ~n27121 & n27185 ;
  assign n27184 = n27121 ^ n27116 ;
  assign n27186 = n27185 ^ n27184 ;
  assign n27187 = x25 & n27186 ;
  assign n27189 = n27188 ^ n27187 ;
  assign n27178 = n27113 ^ n27107 ;
  assign n27179 = n27112 & ~n27178 ;
  assign n27175 = n26413 ^ n26412 ;
  assign n27176 = n27175 ^ n27113 ;
  assign n27177 = n27176 ^ n26509 ;
  assign n27180 = n27179 ^ n27177 ;
  assign n27181 = n27180 ^ n26511 ;
  assign n27174 = n25197 ^ x24 ;
  assign n27182 = n27181 ^ n27174 ;
  assign n27171 = n27115 ^ n27105 ;
  assign n27172 = n27115 ^ n25197 ;
  assign n27173 = n27171 & ~n27172 ;
  assign n27183 = n27182 ^ n27173 ;
  assign n27190 = n27189 ^ n27183 ;
  assign n27162 = n27100 ^ n27051 ;
  assign n27157 = n27099 ^ n27052 ;
  assign n27152 = n27098 ^ n27097 ;
  assign n27143 = n27095 ^ n27054 ;
  assign n27138 = n27094 ^ n27056 ;
  assign n27133 = n27093 ^ n27057 ;
  assign n27128 = n27092 ^ n27058 ;
  assign n27125 = n27091 ^ n27059 ;
  assign n27126 = n26442 ^ n26415 ;
  assign n27127 = ~n27125 & ~n27126 ;
  assign n27129 = n27128 ^ n27127 ;
  assign n27130 = n27128 ^ n26446 ;
  assign n27131 = ~n27129 & n27130 ;
  assign n27132 = n27131 ^ n26446 ;
  assign n27134 = n27133 ^ n27132 ;
  assign n27135 = n27133 ^ n26480 ;
  assign n27136 = ~n27134 & n27135 ;
  assign n27137 = n27136 ^ n26480 ;
  assign n27139 = n27138 ^ n27137 ;
  assign n27140 = n27138 ^ n26522 ;
  assign n27141 = ~n27139 & n27140 ;
  assign n27142 = n27141 ^ n26522 ;
  assign n27144 = n27143 ^ n27142 ;
  assign n27145 = n27143 ^ n26542 ;
  assign n27146 = n27144 & ~n27145 ;
  assign n27147 = n27146 ^ n26542 ;
  assign n27124 = n27096 ^ n27053 ;
  assign n27148 = n27147 ^ n27124 ;
  assign n27149 = n27147 ^ n26562 ;
  assign n27150 = ~n27148 & n27149 ;
  assign n27151 = n27150 ^ n26562 ;
  assign n27153 = n27152 ^ n27151 ;
  assign n27154 = n27152 ^ n26684 ;
  assign n27155 = ~n27153 & n27154 ;
  assign n27156 = n27155 ^ n26684 ;
  assign n27158 = n27157 ^ n27156 ;
  assign n27159 = n27157 ^ n26694 ;
  assign n27160 = ~n27158 & ~n27159 ;
  assign n27161 = n27160 ^ n26694 ;
  assign n27163 = n27162 ^ n27161 ;
  assign n27164 = n27162 ^ n26700 ;
  assign n27165 = ~n27163 & ~n27164 ;
  assign n27166 = n27165 ^ n26700 ;
  assign n27122 = n27121 ^ x25 ;
  assign n27123 = n27122 ^ n27101 ;
  assign n27167 = n27166 ^ n27123 ;
  assign n27168 = n27166 ^ n26706 ;
  assign n27169 = ~n27167 & ~n27168 ;
  assign n27170 = n27169 ^ n26706 ;
  assign n27191 = n27190 ^ n27170 ;
  assign n27192 = n26718 ^ n26712 ;
  assign n27193 = n27192 ^ n26718 ;
  assign n27194 = n27193 ^ n27170 ;
  assign n27195 = n27191 & ~n27194 ;
  assign n27196 = n27195 ^ n27192 ;
  assign n27199 = n26724 ^ n26718 ;
  assign n27197 = n26416 ^ x7 ;
  assign n27198 = n27197 ^ n26724 ;
  assign n27200 = n27199 ^ n27198 ;
  assign n27201 = ~n27196 & n27200 ;
  assign n27202 = n27201 ^ n27199 ;
  assign n27204 = n26730 ^ n26451 ;
  assign n27203 = n26730 ^ n26724 ;
  assign n27205 = n27204 ^ n27203 ;
  assign n27206 = ~n27202 & n27205 ;
  assign n27207 = n27206 ^ n27203 ;
  assign n27210 = n26736 ^ n26730 ;
  assign n27208 = n26492 ^ n26451 ;
  assign n27209 = n27208 ^ n26736 ;
  assign n27211 = n27210 ^ n27209 ;
  assign n27212 = ~n27207 & n27211 ;
  assign n27213 = n27212 ^ n27210 ;
  assign n27216 = n26736 ^ n26656 ;
  assign n27214 = n26534 ^ n26493 ;
  assign n27215 = n27214 ^ n26656 ;
  assign n27217 = n27216 ^ n27215 ;
  assign n27218 = ~n27213 & n27217 ;
  assign n27219 = n27218 ^ n27216 ;
  assign n27220 = ~n26657 & n27219 ;
  assign n27221 = n27220 ^ n26656 ;
  assign n26574 = n26573 ^ n26555 ;
  assign n27222 = n27221 ^ n26574 ;
  assign n27223 = n27061 ^ n27060 ;
  assign n27224 = n27223 ^ n26742 ;
  assign n27225 = n27224 ^ n27223 ;
  assign n27226 = n27225 ^ n26574 ;
  assign n27227 = n27222 & n27226 ;
  assign n27228 = n27227 ^ n27224 ;
  assign n27230 = n26749 ^ n26680 ;
  assign n27229 = n27223 ^ n26680 ;
  assign n27231 = n27230 ^ n27229 ;
  assign n27232 = n27228 & ~n27231 ;
  assign n27233 = n27232 ^ n27230 ;
  assign n27236 = n26771 ^ n26680 ;
  assign n27234 = n27063 ^ n27062 ;
  assign n27235 = n27234 ^ n26771 ;
  assign n27237 = n27236 ^ n27235 ;
  assign n27238 = ~n27233 & ~n27237 ;
  assign n27239 = n27238 ^ n27236 ;
  assign n27243 = n26785 ^ n26771 ;
  assign n27240 = n27065 ^ n27064 ;
  assign n27242 = n27240 ^ n26785 ;
  assign n27244 = n27243 ^ n27242 ;
  assign n27245 = ~n27239 & ~n27244 ;
  assign n27246 = n27245 ^ n27243 ;
  assign n27285 = n26799 ^ n26785 ;
  assign n27247 = n27067 ^ n27066 ;
  assign n27284 = n27247 ^ n26799 ;
  assign n27286 = n27285 ^ n27284 ;
  assign n27287 = n27246 & n27286 ;
  assign n27288 = n27287 ^ n27285 ;
  assign n27291 = n26812 ^ n26799 ;
  assign n27289 = n27069 ^ n27068 ;
  assign n27290 = n27289 ^ n26812 ;
  assign n27292 = n27291 ^ n27290 ;
  assign n27293 = n27288 & n27292 ;
  assign n27294 = n27293 ^ n27291 ;
  assign n27297 = n26823 ^ n26812 ;
  assign n27295 = n27071 ^ n27070 ;
  assign n27296 = n27295 ^ n26823 ;
  assign n27298 = n27297 ^ n27296 ;
  assign n27299 = ~n27294 & ~n27298 ;
  assign n27300 = n27299 ^ n27297 ;
  assign n27282 = n27073 ^ n27072 ;
  assign n27444 = n27300 ^ n27282 ;
  assign n27445 = n27444 ^ n26823 ;
  assign n27446 = n27445 ^ n26000 ;
  assign n27319 = n27295 ^ n27294 ;
  assign n27320 = n27319 ^ n26812 ;
  assign n27321 = n27320 ^ n26805 ;
  assign n27322 = n27321 ^ n25528 ;
  assign n27323 = n27289 ^ n27288 ;
  assign n27324 = n27323 ^ n26799 ;
  assign n27325 = n27324 ^ n26792 ;
  assign n27326 = n27325 ^ n25515 ;
  assign n27248 = n27247 ^ n27246 ;
  assign n27327 = n27248 ^ n26785 ;
  assign n27328 = n27327 ^ n26778 ;
  assign n27329 = n27328 ^ n25383 ;
  assign n27241 = n27240 ^ n27239 ;
  assign n27330 = n27241 ^ n26771 ;
  assign n27331 = n27330 ^ n26764 ;
  assign n27332 = n27331 ^ n25386 ;
  assign n27250 = n27234 ^ n27233 ;
  assign n27333 = n27250 ^ n26680 ;
  assign n27334 = n27333 ^ n26671 ;
  assign n27335 = n27334 ^ n25389 ;
  assign n27408 = n27219 ^ n26575 ;
  assign n27409 = n27408 ^ n26656 ;
  assign n27410 = n27409 ^ n26648 ;
  assign n27336 = n27214 ^ n27213 ;
  assign n27337 = n27336 ^ n26736 ;
  assign n27338 = n27337 ^ n26641 ;
  assign n27339 = n27338 ^ n25393 ;
  assign n27340 = n27208 ^ n27207 ;
  assign n27341 = n27340 ^ n26730 ;
  assign n27342 = n27341 ^ n26633 ;
  assign n27343 = n27342 ^ n25472 ;
  assign n27369 = n27148 ^ n26560 ;
  assign n27364 = n27144 ^ n26538 ;
  assign n27359 = n27139 ^ n26497 ;
  assign n27263 = n27134 ^ n26457 ;
  assign n27253 = n27125 ^ n25923 ;
  assign n27254 = n25924 & n27253 ;
  assign n27255 = n27254 ^ n25401 ;
  assign n27252 = n27129 ^ n26444 ;
  assign n27259 = n27254 ^ n27252 ;
  assign n27260 = ~n27255 & n27259 ;
  assign n27261 = n27260 ^ n25401 ;
  assign n27355 = n27263 ^ n27261 ;
  assign n27356 = n27263 ^ n25407 ;
  assign n27357 = n27355 & n27356 ;
  assign n27358 = n27357 ^ n25407 ;
  assign n27360 = n27359 ^ n27358 ;
  assign n27361 = n27359 ^ n25396 ;
  assign n27362 = n27360 & n27361 ;
  assign n27363 = n27362 ^ n25396 ;
  assign n27365 = n27364 ^ n27363 ;
  assign n27366 = n27364 ^ n25417 ;
  assign n27367 = n27365 & n27366 ;
  assign n27368 = n27367 ^ n25417 ;
  assign n27370 = n27369 ^ n27368 ;
  assign n27371 = n27369 ^ n25423 ;
  assign n27372 = ~n27370 & ~n27371 ;
  assign n27373 = n27372 ^ n25423 ;
  assign n27354 = n27153 ^ n26578 ;
  assign n27374 = n27373 ^ n27354 ;
  assign n27375 = n27373 ^ n25429 ;
  assign n27376 = ~n27374 & n27375 ;
  assign n27377 = n27376 ^ n25429 ;
  assign n27353 = n27158 ^ n26585 ;
  assign n27378 = n27377 ^ n27353 ;
  assign n27379 = n27377 ^ n25435 ;
  assign n27380 = n27378 & ~n27379 ;
  assign n27381 = n27380 ^ n25435 ;
  assign n27352 = n27163 ^ n26593 ;
  assign n27382 = n27381 ^ n27352 ;
  assign n27383 = n27381 ^ n25441 ;
  assign n27384 = n27382 & n27383 ;
  assign n27385 = n27384 ^ n25441 ;
  assign n27351 = n27167 ^ n26601 ;
  assign n27386 = n27385 ^ n27351 ;
  assign n27387 = n27385 ^ n25447 ;
  assign n27388 = ~n27386 & n27387 ;
  assign n27389 = n27388 ^ n25447 ;
  assign n27350 = n27191 ^ n26609 ;
  assign n27390 = n27389 ^ n27350 ;
  assign n27391 = n27389 ^ n25453 ;
  assign n27392 = n27390 & n27391 ;
  assign n27393 = n27392 ^ n25453 ;
  assign n27347 = n27197 ^ n27196 ;
  assign n27348 = n27347 ^ n26718 ;
  assign n27349 = n27348 ^ n26617 ;
  assign n27394 = n27393 ^ n27349 ;
  assign n27395 = n27393 ^ n25459 ;
  assign n27396 = n27394 & n27395 ;
  assign n27397 = n27396 ^ n25459 ;
  assign n27344 = n27202 ^ n26451 ;
  assign n27345 = n27344 ^ n26724 ;
  assign n27346 = n27345 ^ n26625 ;
  assign n27398 = n27397 ^ n27346 ;
  assign n27399 = n27397 ^ n25466 ;
  assign n27400 = ~n27398 & ~n27399 ;
  assign n27401 = n27400 ^ n25466 ;
  assign n27402 = n27401 ^ n27342 ;
  assign n27403 = n27343 & ~n27402 ;
  assign n27404 = n27403 ^ n25472 ;
  assign n27405 = n27404 ^ n27338 ;
  assign n27406 = ~n27339 & n27405 ;
  assign n27407 = n27406 ^ n25393 ;
  assign n27411 = n27410 ^ n27407 ;
  assign n27278 = n26742 ^ n26574 ;
  assign n27279 = n27278 ^ n27221 ;
  assign n27412 = n27279 ^ n26742 ;
  assign n27413 = n27412 ^ n26659 ;
  assign n27414 = n27413 ^ n25480 ;
  assign n27415 = n27414 ^ n27407 ;
  assign n27416 = n27415 ^ n27413 ;
  assign n27417 = n27411 & n27416 ;
  assign n27418 = n27417 ^ n27414 ;
  assign n27419 = n27228 ^ n26673 ;
  assign n27421 = n27419 ^ n25483 ;
  assign n27420 = n27419 ^ n27413 ;
  assign n27422 = n27421 ^ n27420 ;
  assign n27423 = ~n27418 & ~n27422 ;
  assign n27424 = n27423 ^ n27421 ;
  assign n27426 = n27334 ^ n25490 ;
  assign n27425 = n27419 ^ n27334 ;
  assign n27427 = n27426 ^ n27425 ;
  assign n27428 = n27424 & ~n27427 ;
  assign n27429 = n27428 ^ n27426 ;
  assign n27430 = n27335 & n27429 ;
  assign n27431 = n27430 ^ n25389 ;
  assign n27432 = n27431 ^ n27331 ;
  assign n27433 = n27332 & n27432 ;
  assign n27434 = n27433 ^ n25386 ;
  assign n27435 = n27434 ^ n27328 ;
  assign n27436 = ~n27329 & n27435 ;
  assign n27437 = n27436 ^ n25383 ;
  assign n27438 = n27437 ^ n27325 ;
  assign n27439 = n27326 & ~n27438 ;
  assign n27440 = n27439 ^ n25515 ;
  assign n27441 = n27440 ^ n27321 ;
  assign n27442 = n27322 & n27441 ;
  assign n27443 = n27442 ^ n25528 ;
  assign n27447 = n27446 ^ n27443 ;
  assign n27281 = n27075 ^ n27074 ;
  assign n27448 = n27281 ^ n26831 ;
  assign n27283 = n27282 ^ n26823 ;
  assign n27301 = ~n27283 & n27300 ;
  assign n27302 = n27301 ^ n26823 ;
  assign n27449 = n27448 ^ n27302 ;
  assign n27450 = n27449 ^ n26831 ;
  assign n27451 = n27450 ^ n26126 ;
  assign n27452 = n27451 ^ n25539 ;
  assign n27453 = n27452 ^ n27443 ;
  assign n27454 = n27453 ^ n27451 ;
  assign n27455 = ~n27447 & ~n27454 ;
  assign n27456 = n27455 ^ n27452 ;
  assign n27670 = n27456 ^ n25548 ;
  assign n27532 = n27443 ^ n25539 ;
  assign n27533 = n27532 ^ n27446 ;
  assign n27534 = n27533 ^ x112 ;
  assign n27621 = n27418 ^ n25483 ;
  assign n27535 = n27407 ^ n25480 ;
  assign n27536 = n27535 ^ n27410 ;
  assign n27537 = n27536 ^ x104 ;
  assign n27540 = n27399 ^ n27346 ;
  assign n27541 = n27540 ^ x107 ;
  assign n27257 = x103 & ~n27253 ;
  assign n27256 = n27255 ^ n27252 ;
  assign n27258 = n27257 ^ n27256 ;
  assign n27262 = n27261 ^ n25407 ;
  assign n27264 = n27263 ^ n27262 ;
  assign n27265 = n27264 ^ x102 ;
  assign n27266 = n27265 ^ n27256 ;
  assign n27267 = n27266 ^ n27264 ;
  assign n27268 = ~n27258 & n27267 ;
  assign n27269 = n27268 ^ n27265 ;
  assign n27542 = n27358 ^ n25396 ;
  assign n27543 = n27542 ^ n27359 ;
  assign n27545 = n27543 ^ x101 ;
  assign n27544 = n27543 ^ n27264 ;
  assign n27546 = n27545 ^ n27544 ;
  assign n27547 = n27269 & ~n27546 ;
  assign n27548 = n27547 ^ n27545 ;
  assign n27549 = n27363 ^ n25417 ;
  assign n27550 = n27549 ^ n27364 ;
  assign n27552 = n27550 ^ x100 ;
  assign n27551 = n27550 ^ n27543 ;
  assign n27553 = n27552 ^ n27551 ;
  assign n27554 = ~n27548 & n27553 ;
  assign n27555 = n27554 ^ n27552 ;
  assign n27556 = n27368 ^ n25423 ;
  assign n27557 = n27556 ^ n27369 ;
  assign n27559 = n27557 ^ x99 ;
  assign n27558 = n27557 ^ n27550 ;
  assign n27560 = n27559 ^ n27558 ;
  assign n27561 = n27555 & ~n27560 ;
  assign n27562 = n27561 ^ n27559 ;
  assign n27563 = n27375 ^ n27354 ;
  assign n27565 = n27563 ^ x98 ;
  assign n27564 = n27563 ^ n27557 ;
  assign n27566 = n27565 ^ n27564 ;
  assign n27567 = n27562 & ~n27566 ;
  assign n27568 = n27567 ^ n27565 ;
  assign n27569 = n27379 ^ n27353 ;
  assign n27571 = n27569 ^ x97 ;
  assign n27570 = n27569 ^ n27563 ;
  assign n27572 = n27571 ^ n27570 ;
  assign n27573 = n27568 & ~n27572 ;
  assign n27574 = n27573 ^ n27571 ;
  assign n27575 = n27383 ^ n27352 ;
  assign n27577 = n27575 ^ x96 ;
  assign n27576 = n27575 ^ n27569 ;
  assign n27578 = n27577 ^ n27576 ;
  assign n27579 = n27574 & ~n27578 ;
  assign n27580 = n27579 ^ n27577 ;
  assign n27581 = n27387 ^ n27351 ;
  assign n27583 = n27581 ^ x111 ;
  assign n27582 = n27581 ^ n27575 ;
  assign n27584 = n27583 ^ n27582 ;
  assign n27585 = n27580 & ~n27584 ;
  assign n27586 = n27585 ^ n27583 ;
  assign n27587 = n27391 ^ n27350 ;
  assign n27589 = n27587 ^ x110 ;
  assign n27588 = n27587 ^ n27581 ;
  assign n27590 = n27589 ^ n27588 ;
  assign n27591 = ~n27586 & n27590 ;
  assign n27592 = n27591 ^ n27589 ;
  assign n27593 = n27395 ^ n27349 ;
  assign n27595 = n27593 ^ x109 ;
  assign n27594 = n27593 ^ n27587 ;
  assign n27596 = n27595 ^ n27594 ;
  assign n27597 = n27592 & ~n27596 ;
  assign n27598 = n27597 ^ n27595 ;
  assign n27600 = n27540 ^ x108 ;
  assign n27599 = n27593 ^ n27540 ;
  assign n27601 = n27600 ^ n27599 ;
  assign n27602 = n27598 & ~n27601 ;
  assign n27603 = n27602 ^ n27600 ;
  assign n27604 = ~n27541 & n27603 ;
  assign n27605 = n27604 ^ x107 ;
  assign n27538 = n27401 ^ n25472 ;
  assign n27539 = n27538 ^ n27342 ;
  assign n27606 = n27605 ^ n27539 ;
  assign n27607 = n27404 ^ n25393 ;
  assign n27608 = n27607 ^ n27338 ;
  assign n27609 = n27608 ^ x106 ;
  assign n27610 = n27609 ^ n27605 ;
  assign n27611 = n27610 ^ n27608 ;
  assign n27612 = n27606 & n27611 ;
  assign n27613 = n27612 ^ n27609 ;
  assign n27615 = n27536 ^ x105 ;
  assign n27614 = n27608 ^ n27536 ;
  assign n27616 = n27615 ^ n27614 ;
  assign n27617 = ~n27613 & n27616 ;
  assign n27618 = n27617 ^ n27615 ;
  assign n27619 = n27537 & ~n27618 ;
  assign n27620 = n27619 ^ x104 ;
  assign n27622 = n27621 ^ n27620 ;
  assign n27623 = n27424 ^ n25490 ;
  assign n27624 = n27623 ^ x119 ;
  assign n27625 = n27624 ^ n27620 ;
  assign n27626 = n27625 ^ n27623 ;
  assign n27627 = ~n27622 & n27626 ;
  assign n27628 = n27627 ^ n27624 ;
  assign n27629 = n27429 ^ n25389 ;
  assign n27631 = n27629 ^ x118 ;
  assign n27630 = n27629 ^ n27623 ;
  assign n27632 = n27631 ^ n27630 ;
  assign n27633 = n27628 & ~n27632 ;
  assign n27634 = n27633 ^ n27631 ;
  assign n27635 = n27431 ^ n25386 ;
  assign n27636 = n27635 ^ n27331 ;
  assign n27638 = n27636 ^ x117 ;
  assign n27637 = n27636 ^ n27629 ;
  assign n27639 = n27638 ^ n27637 ;
  assign n27640 = ~n27634 & n27639 ;
  assign n27641 = n27640 ^ n27638 ;
  assign n27642 = n27434 ^ n25383 ;
  assign n27643 = n27642 ^ n27328 ;
  assign n27645 = n27643 ^ x116 ;
  assign n27644 = n27643 ^ n27636 ;
  assign n27646 = n27645 ^ n27644 ;
  assign n27647 = n27641 & ~n27646 ;
  assign n27648 = n27647 ^ n27645 ;
  assign n27649 = n27437 ^ n25515 ;
  assign n27650 = n27649 ^ n27325 ;
  assign n27652 = n27650 ^ x115 ;
  assign n27651 = n27650 ^ n27643 ;
  assign n27653 = n27652 ^ n27651 ;
  assign n27654 = n27648 & ~n27653 ;
  assign n27655 = n27654 ^ n27652 ;
  assign n27656 = n27440 ^ n25528 ;
  assign n27657 = n27656 ^ n27321 ;
  assign n27659 = n27657 ^ x114 ;
  assign n27658 = n27657 ^ n27650 ;
  assign n27660 = n27659 ^ n27658 ;
  assign n27661 = ~n27655 & n27660 ;
  assign n27662 = n27661 ^ n27659 ;
  assign n27664 = n27533 ^ x113 ;
  assign n27663 = n27657 ^ n27533 ;
  assign n27665 = n27664 ^ n27663 ;
  assign n27666 = ~n27662 & n27665 ;
  assign n27667 = n27666 ^ n27664 ;
  assign n27668 = n27534 & ~n27667 ;
  assign n27669 = n27668 ^ x112 ;
  assign n27671 = n27670 ^ n27669 ;
  assign n27458 = n26962 ^ n25548 ;
  assign n27303 = n27302 ^ n27281 ;
  assign n27304 = n27077 ^ n27076 ;
  assign n27305 = n27304 ^ n26831 ;
  assign n27306 = n27305 ^ n27281 ;
  assign n27307 = n27306 ^ n27304 ;
  assign n27308 = ~n27303 & n27307 ;
  assign n27309 = n27308 ^ n27305 ;
  assign n27459 = n27458 ^ n27309 ;
  assign n27457 = n27451 ^ n26962 ;
  assign n27460 = n27459 ^ n27457 ;
  assign n27461 = n27460 ^ n27309 ;
  assign n27462 = ~n27456 & ~n27461 ;
  assign n27463 = n27462 ^ n27459 ;
  assign n27672 = n27463 ^ n25561 ;
  assign n27673 = n27672 ^ x127 ;
  assign n27674 = n27673 ^ n27669 ;
  assign n27675 = n27674 ^ n27672 ;
  assign n27676 = n27671 & n27675 ;
  assign n27677 = n27676 ^ n27673 ;
  assign n27318 = n27309 ^ n26290 ;
  assign n27464 = ~n27318 & n27463 ;
  assign n27310 = n27079 ^ n27078 ;
  assign n27312 = n27310 ^ n26963 ;
  assign n27311 = n27310 ^ n27304 ;
  assign n27313 = n27312 ^ n27311 ;
  assign n27314 = n27309 & n27313 ;
  assign n27315 = n27314 ^ n27312 ;
  assign n27316 = n27315 ^ n26976 ;
  assign n27317 = n27316 ^ n25561 ;
  assign n27465 = n27464 ^ n27317 ;
  assign n27678 = n27465 ^ n25574 ;
  assign n27680 = n27678 ^ x126 ;
  assign n27679 = n27678 ^ n27672 ;
  assign n27681 = n27680 ^ n27679 ;
  assign n27682 = ~n27677 & n27681 ;
  assign n27683 = n27682 ^ n27680 ;
  assign n27466 = n27315 ^ n26308 ;
  assign n27467 = ~n27465 & ~n27466 ;
  assign n27468 = n27467 ^ n25574 ;
  assign n27684 = n27468 ^ n25590 ;
  assign n27474 = n27082 ^ n27080 ;
  assign n27470 = n27005 ^ n26983 ;
  assign n27469 = n27310 ^ n27005 ;
  assign n27471 = n27470 ^ n27469 ;
  assign n27472 = ~n27315 & ~n27471 ;
  assign n27473 = n27472 ^ n27470 ;
  assign n27475 = n27474 ^ n27473 ;
  assign n27476 = n27475 ^ n27005 ;
  assign n27477 = n27476 ^ n26328 ;
  assign n27685 = n27684 ^ n27477 ;
  assign n27687 = n27685 ^ x125 ;
  assign n27686 = n27685 ^ n27678 ;
  assign n27688 = n27687 ^ n27686 ;
  assign n27689 = ~n27683 & n27688 ;
  assign n27690 = n27689 ^ n27687 ;
  assign n27478 = n27477 ^ n27468 ;
  assign n27479 = n27477 ^ n25590 ;
  assign n27480 = n27478 & ~n27479 ;
  assign n27481 = n27480 ^ n25590 ;
  assign n27691 = n27481 ^ n25602 ;
  assign n27487 = n27084 ^ n27083 ;
  assign n27483 = n27024 ^ n27005 ;
  assign n27482 = n27474 ^ n27024 ;
  assign n27484 = n27483 ^ n27482 ;
  assign n27485 = n27473 & ~n27484 ;
  assign n27486 = n27485 ^ n27483 ;
  assign n27488 = n27487 ^ n27486 ;
  assign n27489 = n27488 ^ n27024 ;
  assign n27490 = n27489 ^ n26349 ;
  assign n27692 = n27691 ^ n27490 ;
  assign n27694 = n27692 ^ x124 ;
  assign n27693 = n27692 ^ n27685 ;
  assign n27695 = n27694 ^ n27693 ;
  assign n27696 = n27690 & ~n27695 ;
  assign n27697 = n27696 ^ n27694 ;
  assign n27491 = n27490 ^ n27481 ;
  assign n27492 = n27490 ^ n25602 ;
  assign n27493 = n27491 & n27492 ;
  assign n27494 = n27493 ^ n25602 ;
  assign n27698 = n27494 ^ n25614 ;
  assign n27500 = n27086 ^ n27085 ;
  assign n27496 = n27043 ^ n27024 ;
  assign n27495 = n27487 ^ n27043 ;
  assign n27497 = n27496 ^ n27495 ;
  assign n27498 = n27486 & ~n27497 ;
  assign n27499 = n27498 ^ n27496 ;
  assign n27501 = n27500 ^ n27499 ;
  assign n27502 = n27501 ^ n27043 ;
  assign n27503 = n27502 ^ n26430 ;
  assign n27699 = n27698 ^ n27503 ;
  assign n27701 = n27699 ^ x123 ;
  assign n27700 = n27699 ^ n27692 ;
  assign n27702 = n27701 ^ n27700 ;
  assign n27703 = ~n27697 & n27702 ;
  assign n27704 = n27703 ^ n27701 ;
  assign n27504 = n27503 ^ n27494 ;
  assign n27505 = n27503 ^ n25614 ;
  assign n27506 = n27504 & n27505 ;
  assign n27507 = n27506 ^ n25614 ;
  assign n27705 = n27507 ^ n25626 ;
  assign n27513 = n27088 ^ n27087 ;
  assign n27509 = n27114 ^ n27043 ;
  assign n27508 = n27500 ^ n27114 ;
  assign n27510 = n27509 ^ n27508 ;
  assign n27511 = ~n27499 & ~n27510 ;
  assign n27512 = n27511 ^ n27509 ;
  assign n27514 = n27513 ^ n27512 ;
  assign n27515 = n27514 ^ n27114 ;
  assign n27516 = n27515 ^ n27107 ;
  assign n27706 = n27705 ^ n27516 ;
  assign n27708 = n27706 ^ x122 ;
  assign n27707 = n27706 ^ n27699 ;
  assign n27709 = n27708 ^ n27707 ;
  assign n27710 = n27704 & ~n27709 ;
  assign n27711 = n27710 ^ n27708 ;
  assign n27776 = n27711 ^ x121 ;
  assign n27713 = n27562 ^ x98 ;
  assign n27714 = n27555 ^ x99 ;
  assign n27270 = n27269 ^ x101 ;
  assign n27271 = n27253 ^ x103 ;
  assign n27272 = n27257 ^ x102 ;
  assign n27273 = n27272 ^ n27256 ;
  assign n27274 = ~n27271 & n27273 ;
  assign n27715 = n27270 & ~n27274 ;
  assign n27716 = n27548 ^ x100 ;
  assign n27717 = ~n27715 & n27716 ;
  assign n27718 = ~n27714 & n27717 ;
  assign n27719 = ~n27713 & n27718 ;
  assign n27720 = n27568 ^ x97 ;
  assign n27721 = n27719 & ~n27720 ;
  assign n27722 = n27574 ^ x96 ;
  assign n27723 = ~n27721 & n27722 ;
  assign n27724 = n27580 ^ x111 ;
  assign n27725 = ~n27723 & ~n27724 ;
  assign n27726 = n27586 ^ x110 ;
  assign n27727 = n27725 & n27726 ;
  assign n27728 = n27592 ^ x109 ;
  assign n27729 = n27727 & ~n27728 ;
  assign n27730 = n27598 ^ x108 ;
  assign n27731 = n27729 & ~n27730 ;
  assign n27732 = n27603 ^ x107 ;
  assign n27733 = ~n27731 & n27732 ;
  assign n27734 = n27606 ^ x106 ;
  assign n27735 = n27733 & n27734 ;
  assign n27736 = n27613 ^ x105 ;
  assign n27737 = ~n27735 & n27736 ;
  assign n27738 = n27618 ^ x104 ;
  assign n27739 = n27737 & n27738 ;
  assign n27740 = n27620 ^ x119 ;
  assign n27741 = n27740 ^ n27621 ;
  assign n27742 = ~n27739 & ~n27741 ;
  assign n27743 = n27628 ^ x118 ;
  assign n27744 = n27742 & n27743 ;
  assign n27745 = n27634 ^ x117 ;
  assign n27746 = n27744 & ~n27745 ;
  assign n27747 = n27641 ^ x116 ;
  assign n27748 = n27746 & n27747 ;
  assign n27749 = n27648 ^ x115 ;
  assign n27750 = ~n27748 & ~n27749 ;
  assign n27751 = n27655 ^ x114 ;
  assign n27752 = ~n27750 & ~n27751 ;
  assign n27753 = n27662 ^ x113 ;
  assign n27754 = n27752 & ~n27753 ;
  assign n27755 = n27667 ^ x112 ;
  assign n27756 = n27754 & ~n27755 ;
  assign n27757 = n27669 ^ x127 ;
  assign n27758 = n27757 ^ n27670 ;
  assign n27759 = ~n27756 & ~n27758 ;
  assign n27760 = n27677 ^ x126 ;
  assign n27761 = n27759 & n27760 ;
  assign n27762 = n27683 ^ x125 ;
  assign n27763 = ~n27761 & ~n27762 ;
  assign n27764 = n27690 ^ x124 ;
  assign n27765 = ~n27763 & ~n27764 ;
  assign n27766 = n27697 ^ x123 ;
  assign n27767 = ~n27765 & ~n27766 ;
  assign n27768 = n27704 ^ x122 ;
  assign n27769 = ~n27767 & ~n27768 ;
  assign n27777 = n27776 ^ n27769 ;
  assign n27778 = n27777 ^ n27336 ;
  assign n27779 = n27768 ^ n27767 ;
  assign n27780 = n27779 ^ n27340 ;
  assign n27781 = n27766 ^ n27765 ;
  assign n27782 = n27781 ^ n27344 ;
  assign n27783 = n27764 ^ n27763 ;
  assign n27784 = n27783 ^ n27347 ;
  assign n27786 = n27170 ^ n26712 ;
  assign n27787 = n27786 ^ n27190 ;
  assign n27785 = n27762 ^ n27761 ;
  assign n27788 = n27787 ^ n27785 ;
  assign n27791 = n27760 ^ n27759 ;
  assign n27789 = n27168 ^ n27123 ;
  assign n27792 = n27791 ^ n27789 ;
  assign n27795 = n27758 ^ n27756 ;
  assign n27850 = n27795 ^ n27789 ;
  assign n27793 = n27161 ^ n26700 ;
  assign n27794 = n27793 ^ n27162 ;
  assign n27796 = n27795 ^ n27794 ;
  assign n27799 = n27755 ^ n27754 ;
  assign n27847 = n27799 ^ n27794 ;
  assign n27797 = n27156 ^ n26694 ;
  assign n27798 = n27797 ^ n27157 ;
  assign n27800 = n27799 ^ n27798 ;
  assign n27804 = n27753 ^ n27752 ;
  assign n27801 = n27151 ^ n26684 ;
  assign n27802 = n27801 ^ n27152 ;
  assign n27805 = n27804 ^ n27802 ;
  assign n27807 = n27751 ^ n27750 ;
  assign n27842 = n27807 ^ n27802 ;
  assign n27806 = n27149 ^ n27124 ;
  assign n27808 = n27807 ^ n27806 ;
  assign n27812 = n27749 ^ n27748 ;
  assign n27809 = n27142 ^ n26542 ;
  assign n27810 = n27809 ^ n27143 ;
  assign n27813 = n27812 ^ n27810 ;
  assign n27817 = n27747 ^ n27746 ;
  assign n27814 = n27137 ^ n26522 ;
  assign n27815 = n27814 ^ n27138 ;
  assign n27818 = n27817 ^ n27815 ;
  assign n27822 = n27745 ^ n27744 ;
  assign n27819 = n27132 ^ n26480 ;
  assign n27820 = n27819 ^ n27133 ;
  assign n27823 = n27822 ^ n27820 ;
  assign n27827 = n27126 ^ n27125 ;
  assign n27828 = n27741 ^ n27739 ;
  assign n27829 = n27827 & ~n27828 ;
  assign n27824 = n27127 ^ n26446 ;
  assign n27825 = n27824 ^ n27128 ;
  assign n27830 = n27829 ^ n27825 ;
  assign n27831 = n27743 ^ n27742 ;
  assign n27832 = n27831 ^ n27829 ;
  assign n27833 = n27830 & n27832 ;
  assign n27826 = n27825 ^ n27820 ;
  assign n27834 = n27833 ^ n27826 ;
  assign n27835 = n27823 & n27834 ;
  assign n27821 = n27820 ^ n27815 ;
  assign n27836 = n27835 ^ n27821 ;
  assign n27837 = ~n27818 & n27836 ;
  assign n27816 = n27815 ^ n27810 ;
  assign n27838 = n27837 ^ n27816 ;
  assign n27839 = ~n27813 & ~n27838 ;
  assign n27811 = n27810 ^ n27806 ;
  assign n27840 = n27839 ^ n27811 ;
  assign n27841 = ~n27808 & n27840 ;
  assign n27843 = n27842 ^ n27841 ;
  assign n27844 = n27805 & ~n27843 ;
  assign n27803 = n27802 ^ n27798 ;
  assign n27845 = n27844 ^ n27803 ;
  assign n27846 = ~n27800 & n27845 ;
  assign n27848 = n27847 ^ n27846 ;
  assign n27849 = n27796 & ~n27848 ;
  assign n27851 = n27850 ^ n27849 ;
  assign n27852 = ~n27792 & ~n27851 ;
  assign n27790 = n27789 ^ n27787 ;
  assign n27853 = n27852 ^ n27790 ;
  assign n27854 = n27788 & n27853 ;
  assign n27855 = n27854 ^ n27787 ;
  assign n27856 = n27855 ^ n27783 ;
  assign n27857 = n27784 & n27856 ;
  assign n27858 = n27857 ^ n27347 ;
  assign n27859 = n27858 ^ n27781 ;
  assign n27860 = n27782 & n27859 ;
  assign n27861 = n27860 ^ n27344 ;
  assign n27862 = n27861 ^ n27779 ;
  assign n27863 = n27780 & n27862 ;
  assign n27864 = n27863 ^ n27340 ;
  assign n27865 = n27864 ^ n27777 ;
  assign n27866 = n27778 & n27865 ;
  assign n27867 = n27866 ^ n27336 ;
  assign n27869 = n27867 ^ n27408 ;
  assign n27770 = n27769 ^ n27706 ;
  assign n27773 = ~n27711 & ~n27770 ;
  assign n27712 = n27711 ^ n27706 ;
  assign n27771 = n27770 ^ n27712 ;
  assign n27772 = x121 & ~n27771 ;
  assign n27774 = n27773 ^ n27772 ;
  assign n27524 = n27513 ^ n27114 ;
  assign n27525 = ~n27512 & ~n27524 ;
  assign n27522 = n27090 ^ n27089 ;
  assign n27521 = n27513 ^ n27180 ;
  assign n27523 = n27522 ^ n27521 ;
  assign n27526 = n27525 ^ n27523 ;
  assign n27527 = n27526 ^ n27180 ;
  assign n27528 = n27527 ^ n26509 ;
  assign n27529 = n27528 ^ n25637 ;
  assign n27520 = n25626 ^ x120 ;
  assign n27530 = n27529 ^ n27520 ;
  assign n27517 = n27516 ^ n27507 ;
  assign n27518 = n27516 ^ n25626 ;
  assign n27519 = ~n27517 & n27518 ;
  assign n27531 = n27530 ^ n27519 ;
  assign n27775 = n27774 ^ n27531 ;
  assign n28002 = n27869 ^ n27775 ;
  assign n28003 = n28002 ^ n27409 ;
  assign n27912 = n27864 ^ n27336 ;
  assign n27913 = n27912 ^ n27777 ;
  assign n27914 = n27913 ^ n27337 ;
  assign n27915 = n27914 ^ n26641 ;
  assign n27916 = n27861 ^ n27340 ;
  assign n27917 = n27916 ^ n27779 ;
  assign n27918 = n27917 ^ n27341 ;
  assign n27919 = n27918 ^ n26633 ;
  assign n27920 = n27858 ^ n27344 ;
  assign n27921 = n27920 ^ n27781 ;
  assign n27922 = n27921 ^ n27345 ;
  assign n27923 = n27922 ^ n26625 ;
  assign n27924 = n27855 ^ n27347 ;
  assign n27925 = n27924 ^ n27783 ;
  assign n27926 = n27925 ^ n27348 ;
  assign n27927 = n27926 ^ n26617 ;
  assign n27928 = n27853 ^ n27785 ;
  assign n27929 = n27928 ^ n27191 ;
  assign n27930 = n27929 ^ n26609 ;
  assign n27931 = n27851 ^ n27791 ;
  assign n27932 = n27931 ^ n27167 ;
  assign n27933 = n27932 ^ n26601 ;
  assign n27934 = n27848 ^ n27795 ;
  assign n27935 = n27934 ^ n27163 ;
  assign n27936 = n27935 ^ n26593 ;
  assign n27937 = n27845 ^ n27799 ;
  assign n27938 = n27937 ^ n27158 ;
  assign n27939 = n27938 ^ n26585 ;
  assign n27940 = n27843 ^ n27804 ;
  assign n27941 = n27940 ^ n27153 ;
  assign n27942 = n27941 ^ n26578 ;
  assign n27943 = n27840 ^ n27807 ;
  assign n27944 = n27943 ^ n27148 ;
  assign n27945 = n27944 ^ n26560 ;
  assign n27946 = n27838 ^ n27812 ;
  assign n27947 = n27946 ^ n27144 ;
  assign n27948 = n27947 ^ n26538 ;
  assign n27949 = n27828 ^ n27126 ;
  assign n27950 = n26442 & n27949 ;
  assign n27951 = n27950 ^ n26444 ;
  assign n27952 = n27831 ^ n27830 ;
  assign n27953 = n27952 ^ n27129 ;
  assign n27954 = n27953 ^ n27950 ;
  assign n27955 = ~n27951 & n27954 ;
  assign n27956 = n27955 ^ n26444 ;
  assign n27957 = n27956 ^ n26457 ;
  assign n27958 = n27834 ^ n27822 ;
  assign n27959 = n27958 ^ n27134 ;
  assign n27960 = n27959 ^ n27956 ;
  assign n27961 = ~n27957 & n27960 ;
  assign n27962 = n27961 ^ n26457 ;
  assign n27963 = n27962 ^ n26497 ;
  assign n27964 = n27836 ^ n27817 ;
  assign n27965 = n27964 ^ n27139 ;
  assign n27966 = n27965 ^ n27962 ;
  assign n27967 = ~n27963 & n27966 ;
  assign n27968 = n27967 ^ n26497 ;
  assign n27969 = n27968 ^ n27947 ;
  assign n27970 = ~n27948 & n27969 ;
  assign n27971 = n27970 ^ n26538 ;
  assign n27972 = n27971 ^ n27944 ;
  assign n27973 = n27945 & n27972 ;
  assign n27974 = n27973 ^ n26560 ;
  assign n27975 = n27974 ^ n27941 ;
  assign n27976 = n27942 & n27975 ;
  assign n27977 = n27976 ^ n26578 ;
  assign n27978 = n27977 ^ n27938 ;
  assign n27979 = ~n27939 & ~n27978 ;
  assign n27980 = n27979 ^ n26585 ;
  assign n27981 = n27980 ^ n27935 ;
  assign n27982 = ~n27936 & ~n27981 ;
  assign n27983 = n27982 ^ n26593 ;
  assign n27984 = n27983 ^ n27932 ;
  assign n27985 = ~n27933 & ~n27984 ;
  assign n27986 = n27985 ^ n26601 ;
  assign n27987 = n27986 ^ n27929 ;
  assign n27988 = n27930 & ~n27987 ;
  assign n27989 = n27988 ^ n26609 ;
  assign n27990 = n27989 ^ n27926 ;
  assign n27991 = n27927 & ~n27990 ;
  assign n27992 = n27991 ^ n26617 ;
  assign n27993 = n27992 ^ n27922 ;
  assign n27994 = n27923 & n27993 ;
  assign n27995 = n27994 ^ n26625 ;
  assign n27996 = n27995 ^ n27918 ;
  assign n27997 = n27919 & n27996 ;
  assign n27998 = n27997 ^ n26633 ;
  assign n27999 = n27998 ^ n27914 ;
  assign n28000 = n27915 & n27999 ;
  assign n28001 = n28000 ^ n26641 ;
  assign n28004 = n28003 ^ n28001 ;
  assign n27868 = n27867 ^ n27775 ;
  assign n27870 = ~n27868 & n27869 ;
  assign n27871 = n27870 ^ n27408 ;
  assign n28005 = n27871 ^ n27271 ;
  assign n28006 = n28005 ^ n27279 ;
  assign n28007 = n28006 ^ n27412 ;
  assign n28008 = n28007 ^ n26648 ;
  assign n28009 = n28008 ^ n28001 ;
  assign n28010 = n28009 ^ n28007 ;
  assign n28011 = n28004 & n28010 ;
  assign n28012 = n28011 ^ n28008 ;
  assign n28154 = n28012 ^ n26659 ;
  assign n28051 = n28001 ^ n26648 ;
  assign n28052 = n28051 ^ n28003 ;
  assign n28053 = n28052 ^ x200 ;
  assign n28055 = n27828 ^ n26415 ;
  assign n28056 = x199 & n28055 ;
  assign n28054 = n27953 ^ n27951 ;
  assign n28057 = n28056 ^ n28054 ;
  assign n28058 = n27959 ^ n27957 ;
  assign n28059 = n28058 ^ x198 ;
  assign n28060 = n28059 ^ n28054 ;
  assign n28061 = n28060 ^ n28058 ;
  assign n28062 = ~n28057 & n28061 ;
  assign n28063 = n28062 ^ n28059 ;
  assign n28064 = n27965 ^ n27963 ;
  assign n28066 = n28064 ^ x197 ;
  assign n28065 = n28064 ^ n28058 ;
  assign n28067 = n28066 ^ n28065 ;
  assign n28068 = n28063 & ~n28067 ;
  assign n28069 = n28068 ^ n28066 ;
  assign n28070 = n27968 ^ n26538 ;
  assign n28071 = n28070 ^ n27947 ;
  assign n28073 = n28071 ^ x196 ;
  assign n28072 = n28071 ^ n28064 ;
  assign n28074 = n28073 ^ n28072 ;
  assign n28075 = ~n28069 & n28074 ;
  assign n28076 = n28075 ^ n28073 ;
  assign n28077 = n27971 ^ n26560 ;
  assign n28078 = n28077 ^ n27944 ;
  assign n28080 = n28078 ^ x195 ;
  assign n28079 = n28078 ^ n28071 ;
  assign n28081 = n28080 ^ n28079 ;
  assign n28082 = ~n28076 & n28081 ;
  assign n28083 = n28082 ^ n28080 ;
  assign n28084 = n27974 ^ n26578 ;
  assign n28085 = n28084 ^ n27941 ;
  assign n28087 = n28085 ^ x194 ;
  assign n28086 = n28085 ^ n28078 ;
  assign n28088 = n28087 ^ n28086 ;
  assign n28089 = n28083 & ~n28088 ;
  assign n28090 = n28089 ^ n28087 ;
  assign n28091 = n27977 ^ n26585 ;
  assign n28092 = n28091 ^ n27938 ;
  assign n28094 = n28092 ^ x193 ;
  assign n28093 = n28092 ^ n28085 ;
  assign n28095 = n28094 ^ n28093 ;
  assign n28096 = ~n28090 & n28095 ;
  assign n28097 = n28096 ^ n28094 ;
  assign n28098 = n27980 ^ n26593 ;
  assign n28099 = n28098 ^ n27935 ;
  assign n28101 = n28099 ^ x192 ;
  assign n28100 = n28099 ^ n28092 ;
  assign n28102 = n28101 ^ n28100 ;
  assign n28103 = ~n28097 & n28102 ;
  assign n28104 = n28103 ^ n28101 ;
  assign n28105 = n27983 ^ n26601 ;
  assign n28106 = n28105 ^ n27932 ;
  assign n28108 = n28106 ^ x207 ;
  assign n28107 = n28106 ^ n28099 ;
  assign n28109 = n28108 ^ n28107 ;
  assign n28110 = n28104 & ~n28109 ;
  assign n28111 = n28110 ^ n28108 ;
  assign n28112 = n27986 ^ n26609 ;
  assign n28113 = n28112 ^ n27929 ;
  assign n28115 = n28113 ^ x206 ;
  assign n28114 = n28113 ^ n28106 ;
  assign n28116 = n28115 ^ n28114 ;
  assign n28117 = ~n28111 & n28116 ;
  assign n28118 = n28117 ^ n28115 ;
  assign n28119 = n27989 ^ n26617 ;
  assign n28120 = n28119 ^ n27926 ;
  assign n28122 = n28120 ^ x205 ;
  assign n28121 = n28120 ^ n28113 ;
  assign n28123 = n28122 ^ n28121 ;
  assign n28124 = ~n28118 & n28123 ;
  assign n28125 = n28124 ^ n28122 ;
  assign n28126 = n27992 ^ n26625 ;
  assign n28127 = n28126 ^ n27922 ;
  assign n28129 = n28127 ^ x204 ;
  assign n28128 = n28127 ^ n28120 ;
  assign n28130 = n28129 ^ n28128 ;
  assign n28131 = ~n28125 & n28130 ;
  assign n28132 = n28131 ^ n28129 ;
  assign n28133 = n27995 ^ n26633 ;
  assign n28134 = n28133 ^ n27918 ;
  assign n28136 = n28134 ^ x203 ;
  assign n28135 = n28134 ^ n28127 ;
  assign n28137 = n28136 ^ n28135 ;
  assign n28138 = ~n28132 & n28137 ;
  assign n28139 = n28138 ^ n28136 ;
  assign n28140 = n27998 ^ n26641 ;
  assign n28141 = n28140 ^ n27914 ;
  assign n28143 = n28141 ^ x202 ;
  assign n28142 = n28141 ^ n28134 ;
  assign n28144 = n28143 ^ n28142 ;
  assign n28145 = n28139 & ~n28144 ;
  assign n28146 = n28145 ^ n28143 ;
  assign n28148 = n28052 ^ x201 ;
  assign n28147 = n28141 ^ n28052 ;
  assign n28149 = n28148 ^ n28147 ;
  assign n28150 = ~n28146 & n28149 ;
  assign n28151 = n28150 ^ n28148 ;
  assign n28152 = n28053 & ~n28151 ;
  assign n28153 = n28152 ^ x200 ;
  assign n28155 = n28154 ^ n28153 ;
  assign n27876 = n27228 ^ n26749 ;
  assign n27280 = n27279 ^ n27271 ;
  assign n27872 = n27871 ^ n27279 ;
  assign n27873 = n27280 & n27872 ;
  assign n27874 = n27873 ^ n27271 ;
  assign n27277 = n27273 ^ n27271 ;
  assign n27875 = n27874 ^ n27277 ;
  assign n28013 = n27876 ^ n27875 ;
  assign n28014 = n28013 ^ n27228 ;
  assign n28016 = n28014 ^ n26659 ;
  assign n28015 = n28014 ^ n28007 ;
  assign n28017 = n28016 ^ n28015 ;
  assign n28018 = n28012 & n28017 ;
  assign n28019 = n28018 ^ n28016 ;
  assign n28156 = n28019 ^ n26673 ;
  assign n28157 = n28156 ^ x215 ;
  assign n28158 = n28157 ^ n28153 ;
  assign n28159 = n28158 ^ n28156 ;
  assign n28160 = n28155 & n28159 ;
  assign n28161 = n28160 ^ n28157 ;
  assign n27878 = n27874 ^ n27250 ;
  assign n27877 = n27876 ^ n27250 ;
  assign n27879 = n27878 ^ n27877 ;
  assign n27880 = n27875 & n27879 ;
  assign n27881 = n27880 ^ n27877 ;
  assign n27275 = n27274 ^ n27270 ;
  assign n28023 = n27881 ^ n27275 ;
  assign n28024 = n28023 ^ n27333 ;
  assign n28020 = n27875 ^ n26669 ;
  assign n28021 = ~n28019 & n28020 ;
  assign n28022 = n28021 ^ n26673 ;
  assign n28025 = n28024 ^ n28022 ;
  assign n28162 = n28025 ^ n26671 ;
  assign n28164 = n28162 ^ x214 ;
  assign n28163 = n28162 ^ n28156 ;
  assign n28165 = n28164 ^ n28163 ;
  assign n28166 = ~n28161 & n28165 ;
  assign n28167 = n28166 ^ n28164 ;
  assign n28026 = n28022 ^ n26671 ;
  assign n28027 = ~n28025 & ~n28026 ;
  assign n28028 = n28027 ^ n26671 ;
  assign n28168 = n28028 ^ n26764 ;
  assign n27884 = n27716 ^ n27715 ;
  assign n27276 = n27275 ^ n27250 ;
  assign n27882 = n27276 & n27881 ;
  assign n27251 = n27250 ^ n27241 ;
  assign n27883 = n27882 ^ n27251 ;
  assign n27909 = n27884 ^ n27883 ;
  assign n27910 = n27909 ^ n27330 ;
  assign n28169 = n28168 ^ n27910 ;
  assign n28171 = n28169 ^ x213 ;
  assign n28170 = n28169 ^ n28162 ;
  assign n28172 = n28171 ^ n28170 ;
  assign n28173 = n28167 & ~n28172 ;
  assign n28174 = n28173 ^ n28171 ;
  assign n27911 = n27910 ^ n26764 ;
  assign n28029 = n28028 ^ n27910 ;
  assign n28030 = n27911 & n28029 ;
  assign n28031 = n28030 ^ n26764 ;
  assign n28175 = n28031 ^ n26778 ;
  assign n27888 = n27717 ^ n27714 ;
  assign n27885 = n27884 ^ n27241 ;
  assign n27886 = ~n27883 & n27885 ;
  assign n27249 = n27248 ^ n27241 ;
  assign n27887 = n27886 ^ n27249 ;
  assign n27906 = n27888 ^ n27887 ;
  assign n27907 = n27906 ^ n27327 ;
  assign n28176 = n28175 ^ n27907 ;
  assign n28178 = n28176 ^ x212 ;
  assign n28177 = n28176 ^ n28169 ;
  assign n28179 = n28178 ^ n28177 ;
  assign n28180 = n28174 & ~n28179 ;
  assign n28181 = n28180 ^ n28178 ;
  assign n27908 = n27907 ^ n26778 ;
  assign n28032 = n28031 ^ n27907 ;
  assign n28033 = n27908 & n28032 ;
  assign n28034 = n28033 ^ n26778 ;
  assign n28182 = n28034 ^ n26792 ;
  assign n27891 = n27718 ^ n27713 ;
  assign n27892 = n27891 ^ n27248 ;
  assign n27889 = n27888 ^ n27248 ;
  assign n27890 = n27887 & n27889 ;
  assign n27893 = n27892 ^ n27890 ;
  assign n27903 = n27893 ^ n27323 ;
  assign n27904 = n27903 ^ n27324 ;
  assign n28183 = n28182 ^ n27904 ;
  assign n28185 = n28183 ^ x211 ;
  assign n28184 = n28183 ^ n28176 ;
  assign n28186 = n28185 ^ n28184 ;
  assign n28187 = ~n28181 & n28186 ;
  assign n28188 = n28187 ^ n28185 ;
  assign n27905 = n27904 ^ n26792 ;
  assign n28035 = n28034 ^ n27904 ;
  assign n28036 = ~n27905 & ~n28035 ;
  assign n28037 = n28036 ^ n26792 ;
  assign n28189 = n28037 ^ n26805 ;
  assign n27899 = n27720 ^ n27719 ;
  assign n27895 = n27323 ^ n27319 ;
  assign n27894 = n27891 ^ n27319 ;
  assign n27896 = n27895 ^ n27894 ;
  assign n27897 = n27893 & n27896 ;
  assign n27898 = n27897 ^ n27894 ;
  assign n27900 = n27899 ^ n27898 ;
  assign n27901 = n27900 ^ n27320 ;
  assign n28190 = n28189 ^ n27901 ;
  assign n28192 = n28190 ^ x210 ;
  assign n28191 = n28190 ^ n28183 ;
  assign n28193 = n28192 ^ n28191 ;
  assign n28194 = ~n28188 & n28193 ;
  assign n28195 = n28194 ^ n28192 ;
  assign n28045 = n27444 ^ n27319 ;
  assign n28043 = n27899 ^ n27319 ;
  assign n28044 = ~n27898 & ~n28043 ;
  assign n28046 = n28045 ^ n28044 ;
  assign n28042 = n27722 ^ n27721 ;
  assign n28047 = n28046 ^ n28042 ;
  assign n28048 = n28047 ^ n27445 ;
  assign n27902 = n27901 ^ n26805 ;
  assign n28038 = n28037 ^ n27901 ;
  assign n28039 = ~n27902 & ~n28038 ;
  assign n28040 = n28039 ^ n26805 ;
  assign n28041 = n28040 ^ n26000 ;
  assign n28049 = n28048 ^ n28041 ;
  assign n28197 = n28049 ^ x209 ;
  assign n28196 = n28190 ^ n28049 ;
  assign n28198 = n28197 ^ n28196 ;
  assign n28199 = n28195 & ~n28198 ;
  assign n28200 = n28199 ^ n28197 ;
  assign n28286 = n28200 ^ x208 ;
  assign n28239 = n28055 ^ x199 ;
  assign n28240 = n28056 ^ x198 ;
  assign n28241 = n28240 ^ n28054 ;
  assign n28242 = n28239 & n28241 ;
  assign n28243 = n28063 ^ x197 ;
  assign n28244 = ~n28242 & n28243 ;
  assign n28245 = n28069 ^ x196 ;
  assign n28246 = ~n28244 & n28245 ;
  assign n28247 = n28076 ^ x195 ;
  assign n28248 = n28246 & n28247 ;
  assign n28249 = n28083 ^ x194 ;
  assign n28250 = n28248 & ~n28249 ;
  assign n28251 = n28090 ^ x193 ;
  assign n28252 = n28250 & n28251 ;
  assign n28253 = n28097 ^ x192 ;
  assign n28254 = n28252 & n28253 ;
  assign n28255 = n28104 ^ x207 ;
  assign n28256 = ~n28254 & n28255 ;
  assign n28257 = n28111 ^ x206 ;
  assign n28258 = ~n28256 & n28257 ;
  assign n28259 = n28118 ^ x205 ;
  assign n28260 = ~n28258 & ~n28259 ;
  assign n28261 = n28125 ^ x204 ;
  assign n28262 = n28260 & ~n28261 ;
  assign n28263 = n28132 ^ x203 ;
  assign n28264 = n28262 & ~n28263 ;
  assign n28265 = n28139 ^ x202 ;
  assign n28266 = ~n28264 & ~n28265 ;
  assign n28267 = n28146 ^ x201 ;
  assign n28268 = n28266 & n28267 ;
  assign n28269 = n28151 ^ x200 ;
  assign n28270 = n28268 & n28269 ;
  assign n28271 = n28153 ^ x215 ;
  assign n28272 = n28271 ^ n28154 ;
  assign n28273 = n28270 & ~n28272 ;
  assign n28274 = n28161 ^ x214 ;
  assign n28275 = n28273 & n28274 ;
  assign n28276 = n28167 ^ x213 ;
  assign n28277 = n28275 & ~n28276 ;
  assign n28278 = n28174 ^ x212 ;
  assign n28279 = ~n28277 & n28278 ;
  assign n28280 = n28181 ^ x211 ;
  assign n28281 = ~n28279 & n28280 ;
  assign n28282 = n28188 ^ x210 ;
  assign n28283 = n28281 & n28282 ;
  assign n28284 = n28195 ^ x209 ;
  assign n28285 = n28283 & ~n28284 ;
  assign n28294 = n28286 ^ n28285 ;
  assign n28295 = n28294 ^ n27913 ;
  assign n28296 = n28284 ^ n28283 ;
  assign n28297 = n28296 ^ n27917 ;
  assign n28298 = n28282 ^ n28281 ;
  assign n28299 = n28298 ^ n27921 ;
  assign n28300 = n28280 ^ n28279 ;
  assign n28301 = n28300 ^ n27925 ;
  assign n28302 = n28278 ^ n28277 ;
  assign n28303 = n28302 ^ n27928 ;
  assign n28304 = n28276 ^ n28275 ;
  assign n28305 = n28304 ^ n27931 ;
  assign n28306 = n28274 ^ n28273 ;
  assign n28307 = n28306 ^ n27934 ;
  assign n28308 = n28272 ^ n28270 ;
  assign n28309 = n28308 ^ n27937 ;
  assign n28310 = n28269 ^ n28268 ;
  assign n28311 = n28310 ^ n27940 ;
  assign n28312 = n28267 ^ n28266 ;
  assign n28313 = n28312 ^ n27943 ;
  assign n28314 = n28265 ^ n28264 ;
  assign n28315 = n28314 ^ n27946 ;
  assign n28316 = n28263 ^ n28262 ;
  assign n28317 = n28316 ^ n27964 ;
  assign n28318 = n28261 ^ n28260 ;
  assign n28319 = n28318 ^ n27958 ;
  assign n28320 = n27949 ^ n27125 ;
  assign n28321 = n28257 ^ n28256 ;
  assign n28322 = ~n28320 & ~n28321 ;
  assign n28323 = n28322 ^ n27952 ;
  assign n28324 = n28259 ^ n28258 ;
  assign n28325 = n28324 ^ n28322 ;
  assign n28326 = ~n28323 & n28325 ;
  assign n28327 = n28326 ^ n27952 ;
  assign n28328 = n28327 ^ n28318 ;
  assign n28329 = n28319 & n28328 ;
  assign n28330 = n28329 ^ n27958 ;
  assign n28331 = n28330 ^ n28316 ;
  assign n28332 = ~n28317 & ~n28331 ;
  assign n28333 = n28332 ^ n27964 ;
  assign n28334 = n28333 ^ n28314 ;
  assign n28335 = ~n28315 & n28334 ;
  assign n28336 = n28335 ^ n27946 ;
  assign n28337 = n28336 ^ n28312 ;
  assign n28338 = n28313 & n28337 ;
  assign n28339 = n28338 ^ n27943 ;
  assign n28340 = n28339 ^ n28310 ;
  assign n28341 = ~n28311 & ~n28340 ;
  assign n28342 = n28341 ^ n27940 ;
  assign n28343 = n28342 ^ n28308 ;
  assign n28344 = n28309 & ~n28343 ;
  assign n28345 = n28344 ^ n27937 ;
  assign n28346 = n28345 ^ n28306 ;
  assign n28347 = n28307 & n28346 ;
  assign n28348 = n28347 ^ n27934 ;
  assign n28349 = n28348 ^ n28304 ;
  assign n28350 = n28305 & n28349 ;
  assign n28351 = n28350 ^ n27931 ;
  assign n28352 = n28351 ^ n28302 ;
  assign n28353 = ~n28303 & n28352 ;
  assign n28354 = n28353 ^ n27928 ;
  assign n28355 = n28354 ^ n28300 ;
  assign n28356 = n28301 & ~n28355 ;
  assign n28357 = n28356 ^ n27925 ;
  assign n28358 = n28357 ^ n28298 ;
  assign n28359 = n28299 & n28358 ;
  assign n28360 = n28359 ^ n27921 ;
  assign n28361 = n28360 ^ n28296 ;
  assign n28362 = n28297 & n28361 ;
  assign n28363 = n28362 ^ n27917 ;
  assign n28364 = n28363 ^ n28294 ;
  assign n28365 = n28295 & n28364 ;
  assign n28366 = n28365 ^ n27913 ;
  assign n28050 = n28049 ^ x208 ;
  assign n28201 = ~n28050 & n28200 ;
  assign n28202 = n28201 ^ x208 ;
  assign n28288 = n28202 ^ x223 ;
  assign n28203 = n28048 ^ n28040 ;
  assign n28209 = n27724 ^ n27723 ;
  assign n28204 = n27449 ^ n27444 ;
  assign n28205 = n28204 ^ n27449 ;
  assign n28206 = n28205 ^ n28042 ;
  assign n28207 = ~n28046 & ~n28206 ;
  assign n28208 = n28207 ^ n28204 ;
  assign n28210 = n28209 ^ n28208 ;
  assign n28211 = n28210 ^ n27450 ;
  assign n28212 = n28211 ^ n26000 ;
  assign n28213 = n28212 ^ n28040 ;
  assign n28214 = n28213 ^ n28211 ;
  assign n28215 = n28203 & ~n28214 ;
  assign n28216 = n28215 ^ n28212 ;
  assign n28217 = n28216 ^ n26126 ;
  assign n28289 = n28288 ^ n28217 ;
  assign n28287 = ~n28285 & n28286 ;
  assign n28292 = n28289 ^ n28287 ;
  assign n28367 = n28366 ^ n28292 ;
  assign n28782 = n28367 ^ n27408 ;
  assign n28580 = n28364 ^ n27336 ;
  assign n28778 = n28580 ^ n26736 ;
  assign n28568 = n28361 ^ n27340 ;
  assign n28575 = n28568 ^ n26730 ;
  assign n28556 = n28358 ^ n27344 ;
  assign n28563 = n28556 ^ n26724 ;
  assign n28544 = n28355 ^ n27347 ;
  assign n28551 = n28544 ^ n26718 ;
  assign n28532 = n28352 ^ n27787 ;
  assign n28539 = n28532 ^ n26712 ;
  assign n28520 = n28349 ^ n27789 ;
  assign n28527 = n28520 ^ n26706 ;
  assign n28508 = n28346 ^ n27794 ;
  assign n28515 = n28508 ^ n26700 ;
  assign n28496 = n28343 ^ n27798 ;
  assign n28503 = n28496 ^ n26694 ;
  assign n28484 = n28340 ^ n27802 ;
  assign n28491 = n28484 ^ n26684 ;
  assign n28472 = n28337 ^ n27806 ;
  assign n28479 = n28472 ^ n26562 ;
  assign n28460 = n28334 ^ n27810 ;
  assign n28467 = n28460 ^ n26542 ;
  assign n28448 = n28331 ^ n27815 ;
  assign n28455 = n28448 ^ n26522 ;
  assign n28436 = n28328 ^ n27820 ;
  assign n28443 = n28436 ^ n26480 ;
  assign n28426 = n28321 ^ n27125 ;
  assign n28427 = ~n27126 & ~n28426 ;
  assign n28428 = n28427 ^ n26446 ;
  assign n28425 = n28325 ^ n27825 ;
  assign n28432 = n28427 ^ n28425 ;
  assign n28433 = n28428 & n28432 ;
  assign n28434 = n28433 ^ n26446 ;
  assign n28444 = n28436 ^ n28434 ;
  assign n28445 = ~n28443 & n28444 ;
  assign n28446 = n28445 ^ n26480 ;
  assign n28456 = n28448 ^ n28446 ;
  assign n28457 = n28455 & ~n28456 ;
  assign n28458 = n28457 ^ n26522 ;
  assign n28468 = n28460 ^ n28458 ;
  assign n28469 = n28467 & ~n28468 ;
  assign n28470 = n28469 ^ n26542 ;
  assign n28480 = n28472 ^ n28470 ;
  assign n28481 = ~n28479 & n28480 ;
  assign n28482 = n28481 ^ n26562 ;
  assign n28492 = n28484 ^ n28482 ;
  assign n28493 = n28491 & ~n28492 ;
  assign n28494 = n28493 ^ n26684 ;
  assign n28504 = n28496 ^ n28494 ;
  assign n28505 = n28503 & n28504 ;
  assign n28506 = n28505 ^ n26694 ;
  assign n28516 = n28508 ^ n28506 ;
  assign n28517 = ~n28515 & ~n28516 ;
  assign n28518 = n28517 ^ n26700 ;
  assign n28528 = n28520 ^ n28518 ;
  assign n28529 = ~n28527 & ~n28528 ;
  assign n28530 = n28529 ^ n26706 ;
  assign n28540 = n28532 ^ n28530 ;
  assign n28541 = n28539 & n28540 ;
  assign n28542 = n28541 ^ n26712 ;
  assign n28552 = n28544 ^ n28542 ;
  assign n28553 = ~n28551 & ~n28552 ;
  assign n28554 = n28553 ^ n26718 ;
  assign n28564 = n28556 ^ n28554 ;
  assign n28565 = n28563 & n28564 ;
  assign n28566 = n28565 ^ n26724 ;
  assign n28576 = n28568 ^ n28566 ;
  assign n28577 = n28575 & n28576 ;
  assign n28578 = n28577 ^ n26730 ;
  assign n28779 = n28580 ^ n28578 ;
  assign n28780 = n28778 & n28779 ;
  assign n28781 = n28780 ^ n26736 ;
  assign n28783 = n28782 ^ n28781 ;
  assign n28293 = n28292 ^ n28002 ;
  assign n28368 = ~n28293 & ~n28367 ;
  assign n28369 = n28368 ^ n28002 ;
  assign n28290 = ~n28287 & ~n28289 ;
  assign n28218 = n28217 ^ n28202 ;
  assign n28224 = n27309 ^ n26963 ;
  assign n28220 = n28209 ^ n27449 ;
  assign n28221 = ~n28208 & n28220 ;
  assign n28222 = n28221 ^ n27449 ;
  assign n28219 = n27726 ^ n27725 ;
  assign n28223 = n28222 ^ n28219 ;
  assign n28225 = n28224 ^ n28223 ;
  assign n28226 = n28225 ^ n27309 ;
  assign n28228 = n28226 ^ n26126 ;
  assign n28227 = n28226 ^ n28211 ;
  assign n28229 = n28228 ^ n28227 ;
  assign n28230 = n28216 & ~n28229 ;
  assign n28231 = n28230 ^ n28228 ;
  assign n28232 = n28231 ^ n26962 ;
  assign n28233 = n28232 ^ x223 ;
  assign n28234 = n28233 ^ n28202 ;
  assign n28235 = n28234 ^ n28232 ;
  assign n28236 = n28218 & n28235 ;
  assign n28237 = n28236 ^ n28233 ;
  assign n28238 = n28237 ^ x222 ;
  assign n28291 = n28290 ^ n28238 ;
  assign n28370 = n28369 ^ n28291 ;
  assign n28784 = n28370 ^ n27279 ;
  assign n28785 = n28784 ^ n26656 ;
  assign n28786 = n28785 ^ n28781 ;
  assign n28787 = n28786 ^ n28784 ;
  assign n28788 = n28783 & n28787 ;
  assign n28789 = n28788 ^ n28785 ;
  assign n28897 = n28789 ^ n26742 ;
  assign n28887 = n28781 ^ n26656 ;
  assign n28888 = n28887 ^ n28782 ;
  assign n28889 = n28888 ^ x296 ;
  assign n28430 = x295 & n28426 ;
  assign n28429 = n28428 ^ n28425 ;
  assign n28431 = n28430 ^ n28429 ;
  assign n28435 = n28434 ^ n26480 ;
  assign n28437 = n28436 ^ n28435 ;
  assign n28438 = n28437 ^ x294 ;
  assign n28439 = n28438 ^ n28429 ;
  assign n28440 = n28439 ^ n28437 ;
  assign n28441 = n28431 & ~n28440 ;
  assign n28442 = n28441 ^ n28438 ;
  assign n28447 = n28446 ^ n26522 ;
  assign n28449 = n28448 ^ n28447 ;
  assign n28451 = n28449 ^ x293 ;
  assign n28450 = n28449 ^ n28437 ;
  assign n28452 = n28451 ^ n28450 ;
  assign n28453 = n28442 & ~n28452 ;
  assign n28454 = n28453 ^ n28451 ;
  assign n28459 = n28458 ^ n26542 ;
  assign n28461 = n28460 ^ n28459 ;
  assign n28463 = n28461 ^ x292 ;
  assign n28462 = n28461 ^ n28449 ;
  assign n28464 = n28463 ^ n28462 ;
  assign n28465 = ~n28454 & n28464 ;
  assign n28466 = n28465 ^ n28463 ;
  assign n28471 = n28470 ^ n26562 ;
  assign n28473 = n28472 ^ n28471 ;
  assign n28475 = n28473 ^ x291 ;
  assign n28474 = n28473 ^ n28461 ;
  assign n28476 = n28475 ^ n28474 ;
  assign n28477 = ~n28466 & n28476 ;
  assign n28478 = n28477 ^ n28475 ;
  assign n28483 = n28482 ^ n26684 ;
  assign n28485 = n28484 ^ n28483 ;
  assign n28487 = n28485 ^ x290 ;
  assign n28486 = n28485 ^ n28473 ;
  assign n28488 = n28487 ^ n28486 ;
  assign n28489 = n28478 & ~n28488 ;
  assign n28490 = n28489 ^ n28487 ;
  assign n28495 = n28494 ^ n26694 ;
  assign n28497 = n28496 ^ n28495 ;
  assign n28499 = n28497 ^ x289 ;
  assign n28498 = n28497 ^ n28485 ;
  assign n28500 = n28499 ^ n28498 ;
  assign n28501 = ~n28490 & n28500 ;
  assign n28502 = n28501 ^ n28499 ;
  assign n28507 = n28506 ^ n26700 ;
  assign n28509 = n28508 ^ n28507 ;
  assign n28511 = n28509 ^ x288 ;
  assign n28510 = n28509 ^ n28497 ;
  assign n28512 = n28511 ^ n28510 ;
  assign n28513 = ~n28502 & n28512 ;
  assign n28514 = n28513 ^ n28511 ;
  assign n28519 = n28518 ^ n26706 ;
  assign n28521 = n28520 ^ n28519 ;
  assign n28523 = n28521 ^ x303 ;
  assign n28522 = n28521 ^ n28509 ;
  assign n28524 = n28523 ^ n28522 ;
  assign n28525 = ~n28514 & n28524 ;
  assign n28526 = n28525 ^ n28523 ;
  assign n28531 = n28530 ^ n26712 ;
  assign n28533 = n28532 ^ n28531 ;
  assign n28535 = n28533 ^ x302 ;
  assign n28534 = n28533 ^ n28521 ;
  assign n28536 = n28535 ^ n28534 ;
  assign n28537 = n28526 & ~n28536 ;
  assign n28538 = n28537 ^ n28535 ;
  assign n28543 = n28542 ^ n26718 ;
  assign n28545 = n28544 ^ n28543 ;
  assign n28547 = n28545 ^ x301 ;
  assign n28546 = n28545 ^ n28533 ;
  assign n28548 = n28547 ^ n28546 ;
  assign n28549 = n28538 & ~n28548 ;
  assign n28550 = n28549 ^ n28547 ;
  assign n28555 = n28554 ^ n26724 ;
  assign n28557 = n28556 ^ n28555 ;
  assign n28559 = n28557 ^ x300 ;
  assign n28558 = n28557 ^ n28545 ;
  assign n28560 = n28559 ^ n28558 ;
  assign n28561 = n28550 & ~n28560 ;
  assign n28562 = n28561 ^ n28559 ;
  assign n28567 = n28566 ^ n26730 ;
  assign n28569 = n28568 ^ n28567 ;
  assign n28571 = n28569 ^ x299 ;
  assign n28570 = n28569 ^ n28557 ;
  assign n28572 = n28571 ^ n28570 ;
  assign n28573 = n28562 & ~n28572 ;
  assign n28574 = n28573 ^ n28571 ;
  assign n28579 = n28578 ^ n26736 ;
  assign n28581 = n28580 ^ n28579 ;
  assign n28583 = n28581 ^ x298 ;
  assign n28582 = n28581 ^ n28569 ;
  assign n28584 = n28583 ^ n28582 ;
  assign n28585 = ~n28574 & n28584 ;
  assign n28586 = n28585 ^ n28583 ;
  assign n28891 = n28888 ^ x297 ;
  assign n28890 = n28888 ^ n28581 ;
  assign n28892 = n28891 ^ n28890 ;
  assign n28893 = n28586 & ~n28892 ;
  assign n28894 = n28893 ^ n28891 ;
  assign n28895 = ~n28889 & n28894 ;
  assign n28896 = n28895 ^ x296 ;
  assign n28898 = n28897 ^ n28896 ;
  assign n28792 = n27876 ^ n26742 ;
  assign n28392 = n28238 & n28290 ;
  assign n28377 = n27728 ^ n27727 ;
  assign n28371 = n27315 ^ n26983 ;
  assign n28372 = n28371 ^ n28224 ;
  assign n28373 = n28372 ^ n28219 ;
  assign n28374 = n28373 ^ n28371 ;
  assign n28375 = ~n28223 & n28374 ;
  assign n28376 = n28375 ^ n28372 ;
  assign n28378 = n28377 ^ n28376 ;
  assign n28379 = n28378 ^ n27315 ;
  assign n28381 = n28379 ^ n26962 ;
  assign n28380 = n28379 ^ n28226 ;
  assign n28382 = n28381 ^ n28380 ;
  assign n28383 = n28231 & n28382 ;
  assign n28384 = n28383 ^ n28381 ;
  assign n28385 = n28384 ^ n26976 ;
  assign n28387 = n28385 ^ x222 ;
  assign n28386 = n28385 ^ n28232 ;
  assign n28388 = n28387 ^ n28386 ;
  assign n28389 = ~n28237 & n28388 ;
  assign n28390 = n28389 ^ n28387 ;
  assign n28391 = n28390 ^ x221 ;
  assign n28393 = n28392 ^ n28391 ;
  assign n28394 = n28393 ^ n28006 ;
  assign n28395 = n28394 ^ n28291 ;
  assign n28396 = n28395 ^ n28393 ;
  assign n28397 = n28370 & ~n28396 ;
  assign n28398 = n28397 ^ n28394 ;
  assign n28793 = n28792 ^ n28398 ;
  assign n28790 = n28784 ^ n27876 ;
  assign n28791 = n28790 ^ n28398 ;
  assign n28794 = n28793 ^ n28791 ;
  assign n28795 = n28789 & n28794 ;
  assign n28796 = n28795 ^ n28793 ;
  assign n28899 = n28796 ^ n26749 ;
  assign n28900 = n28899 ^ x311 ;
  assign n28901 = n28900 ^ n28896 ;
  assign n28902 = n28901 ^ n28899 ;
  assign n28903 = ~n28898 & n28902 ;
  assign n28904 = n28903 ^ n28900 ;
  assign n28777 = n28398 ^ n27228 ;
  assign n28797 = n28777 & ~n28796 ;
  assign n28418 = n28391 & ~n28392 ;
  assign n28403 = n27730 ^ n27729 ;
  assign n28405 = n28403 ^ n28371 ;
  assign n28404 = n28403 ^ n28377 ;
  assign n28406 = n28405 ^ n28404 ;
  assign n28407 = n28376 & ~n28406 ;
  assign n28408 = n28407 ^ n28405 ;
  assign n28409 = n28408 ^ n27475 ;
  assign n28410 = n28409 ^ n27476 ;
  assign n28399 = n28379 ^ n26976 ;
  assign n28400 = ~n28384 & n28399 ;
  assign n28401 = n28400 ^ n26976 ;
  assign n28402 = n28401 ^ n26328 ;
  assign n28411 = n28410 ^ n28402 ;
  assign n28413 = n28411 ^ x221 ;
  assign n28412 = n28411 ^ n28385 ;
  assign n28414 = n28413 ^ n28412 ;
  assign n28415 = n28390 & ~n28414 ;
  assign n28416 = n28415 ^ n28413 ;
  assign n28417 = n28416 ^ x220 ;
  assign n28419 = n28418 ^ n28417 ;
  assign n28421 = n28419 ^ n28013 ;
  assign n28420 = n28419 ^ n28393 ;
  assign n28422 = n28421 ^ n28420 ;
  assign n28423 = n28398 & ~n28422 ;
  assign n28424 = n28423 ^ n28421 ;
  assign n28775 = n28424 ^ n27250 ;
  assign n28776 = n28775 ^ n26749 ;
  assign n28798 = n28797 ^ n28776 ;
  assign n28905 = n28798 ^ n26680 ;
  assign n28907 = n28905 ^ x310 ;
  assign n28906 = n28905 ^ n28899 ;
  assign n28908 = n28907 ^ n28906 ;
  assign n28909 = n28904 & ~n28908 ;
  assign n28910 = n28909 ^ n28907 ;
  assign n28701 = n28419 ^ n28023 ;
  assign n28702 = ~n28424 & ~n28701 ;
  assign n28703 = n28702 ^ n28023 ;
  assign n28642 = n27732 ^ n27731 ;
  assign n28638 = n27488 ^ n27475 ;
  assign n28637 = n28403 ^ n27488 ;
  assign n28639 = n28638 ^ n28637 ;
  assign n28640 = n28408 & n28639 ;
  assign n28641 = n28640 ^ n28638 ;
  assign n28643 = n28642 ^ n28641 ;
  assign n28644 = n28643 ^ n27489 ;
  assign n28632 = n28410 ^ n28401 ;
  assign n28633 = n28410 ^ n26328 ;
  assign n28634 = ~n28632 & ~n28633 ;
  assign n28635 = n28634 ^ n26328 ;
  assign n28636 = n28635 ^ n26349 ;
  assign n28645 = n28644 ^ n28636 ;
  assign n28647 = n28645 ^ x220 ;
  assign n28646 = n28645 ^ n28411 ;
  assign n28648 = n28647 ^ n28646 ;
  assign n28649 = ~n28416 & n28648 ;
  assign n28650 = n28649 ^ n28647 ;
  assign n28691 = n28650 ^ x219 ;
  assign n28690 = n28417 & ~n28418 ;
  assign n28699 = n28691 ^ n28690 ;
  assign n28704 = n28703 ^ n28699 ;
  assign n28803 = n28704 ^ n27241 ;
  assign n28799 = n28775 ^ n26680 ;
  assign n28800 = n28798 & n28799 ;
  assign n28801 = n28800 ^ n26680 ;
  assign n28802 = n28801 ^ n26771 ;
  assign n28911 = n28803 ^ n28802 ;
  assign n28913 = n28911 ^ x309 ;
  assign n28912 = n28911 ^ n28905 ;
  assign n28914 = n28913 ^ n28912 ;
  assign n28915 = n28910 & ~n28914 ;
  assign n28916 = n28915 ^ n28913 ;
  assign n28804 = n28803 ^ n28801 ;
  assign n28805 = ~n28802 & ~n28804 ;
  assign n28806 = n28805 ^ n26771 ;
  assign n28917 = n28806 ^ n26785 ;
  assign n28700 = n28699 ^ n27909 ;
  assign n28705 = ~n28700 & n28704 ;
  assign n28706 = n28705 ^ n27909 ;
  assign n28661 = n27734 ^ n27733 ;
  assign n28657 = n27501 ^ n27488 ;
  assign n28656 = n28642 ^ n27501 ;
  assign n28658 = n28657 ^ n28656 ;
  assign n28659 = n28641 & ~n28658 ;
  assign n28660 = n28659 ^ n28657 ;
  assign n28662 = n28661 ^ n28660 ;
  assign n28663 = n28662 ^ n27502 ;
  assign n28651 = n28644 ^ n28635 ;
  assign n28652 = n28644 ^ n26349 ;
  assign n28653 = n28651 & ~n28652 ;
  assign n28654 = n28653 ^ n26349 ;
  assign n28655 = n28654 ^ n26430 ;
  assign n28664 = n28663 ^ n28655 ;
  assign n28666 = n28664 ^ x219 ;
  assign n28665 = n28664 ^ n28645 ;
  assign n28667 = n28666 ^ n28665 ;
  assign n28668 = n28650 & ~n28667 ;
  assign n28669 = n28668 ^ n28666 ;
  assign n28693 = n28669 ^ x218 ;
  assign n28692 = n28690 & ~n28691 ;
  assign n28697 = n28693 ^ n28692 ;
  assign n28707 = n28706 ^ n28697 ;
  assign n28773 = n28707 ^ n27248 ;
  assign n28918 = n28917 ^ n28773 ;
  assign n28920 = n28918 ^ x308 ;
  assign n28919 = n28918 ^ n28911 ;
  assign n28921 = n28920 ^ n28919 ;
  assign n28922 = n28916 & ~n28921 ;
  assign n28923 = n28922 ^ n28920 ;
  assign n28774 = n28773 ^ n26785 ;
  assign n28807 = n28806 ^ n28773 ;
  assign n28808 = ~n28774 & n28807 ;
  assign n28809 = n28808 ^ n26785 ;
  assign n28924 = n28809 ^ n26799 ;
  assign n28698 = n28697 ^ n27906 ;
  assign n28708 = n28698 & n28707 ;
  assign n28709 = n28708 ^ n27906 ;
  assign n28694 = n28692 & ~n28693 ;
  assign n28680 = n27736 ^ n27735 ;
  assign n28676 = n27514 ^ n27501 ;
  assign n28675 = n28661 ^ n27514 ;
  assign n28677 = n28676 ^ n28675 ;
  assign n28678 = n28660 & n28677 ;
  assign n28679 = n28678 ^ n28676 ;
  assign n28681 = n28680 ^ n28679 ;
  assign n28682 = n28681 ^ n27515 ;
  assign n28670 = n28663 ^ n28654 ;
  assign n28671 = n28663 ^ n26430 ;
  assign n28672 = n28670 & ~n28671 ;
  assign n28673 = n28672 ^ n26430 ;
  assign n28674 = n28673 ^ n27107 ;
  assign n28683 = n28682 ^ n28674 ;
  assign n28685 = n28683 ^ x218 ;
  assign n28684 = n28683 ^ n28664 ;
  assign n28686 = n28685 ^ n28684 ;
  assign n28687 = n28669 & ~n28686 ;
  assign n28688 = n28687 ^ n28685 ;
  assign n28689 = n28688 ^ x217 ;
  assign n28695 = n28694 ^ n28689 ;
  assign n28710 = n28709 ^ n28695 ;
  assign n28771 = n28710 ^ n27323 ;
  assign n28925 = n28924 ^ n28771 ;
  assign n28927 = n28925 ^ x307 ;
  assign n28926 = n28925 ^ n28918 ;
  assign n28928 = n28927 ^ n28926 ;
  assign n28929 = ~n28923 & n28928 ;
  assign n28930 = n28929 ^ n28927 ;
  assign n28772 = n28771 ^ n26799 ;
  assign n28810 = n28809 ^ n28771 ;
  assign n28811 = ~n28772 & n28810 ;
  assign n28812 = n28811 ^ n26799 ;
  assign n28931 = n28812 ^ n26812 ;
  assign n28727 = n28694 ^ n28683 ;
  assign n28730 = ~n28688 & ~n28727 ;
  assign n28726 = n28688 ^ n28683 ;
  assign n28728 = n28727 ^ n28726 ;
  assign n28729 = ~x217 & n28728 ;
  assign n28731 = n28730 ^ n28729 ;
  assign n28720 = n28680 ^ n27514 ;
  assign n28721 = n28679 & ~n28720 ;
  assign n28718 = n27738 ^ n27737 ;
  assign n28717 = n28680 ^ n27526 ;
  assign n28719 = n28718 ^ n28717 ;
  assign n28722 = n28721 ^ n28719 ;
  assign n28723 = n28722 ^ n27528 ;
  assign n28716 = n27107 ^ x216 ;
  assign n28724 = n28723 ^ n28716 ;
  assign n28713 = n28682 ^ n28673 ;
  assign n28714 = n28682 ^ n27107 ;
  assign n28715 = n28713 & n28714 ;
  assign n28725 = n28724 ^ n28715 ;
  assign n28732 = n28731 ^ n28725 ;
  assign n28696 = n28695 ^ n27903 ;
  assign n28711 = ~n28696 & n28710 ;
  assign n28712 = n28711 ^ n27903 ;
  assign n28733 = n28732 ^ n28712 ;
  assign n28769 = n28733 ^ n27319 ;
  assign n28932 = n28931 ^ n28769 ;
  assign n28934 = n28932 ^ x306 ;
  assign n28933 = n28932 ^ n28925 ;
  assign n28935 = n28934 ^ n28933 ;
  assign n28936 = ~n28930 & n28935 ;
  assign n28937 = n28936 ^ n28934 ;
  assign n28770 = n28769 ^ n26812 ;
  assign n28813 = n28812 ^ n28769 ;
  assign n28814 = n28770 & n28813 ;
  assign n28815 = n28814 ^ n26812 ;
  assign n28884 = n28815 ^ n26823 ;
  assign n28734 = n28732 ^ n27900 ;
  assign n28735 = ~n28733 & ~n28734 ;
  assign n28736 = n28735 ^ n27900 ;
  assign n28631 = n28239 ^ n28047 ;
  assign n28766 = n28736 ^ n28631 ;
  assign n28767 = n28766 ^ n28047 ;
  assign n28768 = n28767 ^ n27444 ;
  assign n28885 = n28884 ^ n28768 ;
  assign n28939 = n28885 ^ x305 ;
  assign n28938 = n28932 ^ n28885 ;
  assign n28940 = n28939 ^ n28938 ;
  assign n28941 = n28937 & ~n28940 ;
  assign n28942 = n28941 ^ n28939 ;
  assign n29005 = n28942 ^ x304 ;
  assign n28987 = n28916 ^ x308 ;
  assign n28587 = n28586 ^ x297 ;
  assign n28588 = n28426 ^ x295 ;
  assign n28589 = n28430 ^ x294 ;
  assign n28590 = n28589 ^ n28429 ;
  assign n28591 = n28588 & ~n28590 ;
  assign n28592 = n28442 ^ x293 ;
  assign n28593 = n28591 & ~n28592 ;
  assign n28594 = n28454 ^ x292 ;
  assign n28595 = ~n28593 & ~n28594 ;
  assign n28596 = n28466 ^ x291 ;
  assign n28597 = n28595 & ~n28596 ;
  assign n28598 = n28478 ^ x290 ;
  assign n28599 = n28597 & n28598 ;
  assign n28600 = n28490 ^ x289 ;
  assign n28601 = ~n28599 & n28600 ;
  assign n28602 = n28502 ^ x288 ;
  assign n28603 = n28601 & n28602 ;
  assign n28604 = n28514 ^ x303 ;
  assign n28605 = n28603 & n28604 ;
  assign n28606 = n28526 ^ x302 ;
  assign n28607 = n28605 & ~n28606 ;
  assign n28608 = n28538 ^ x301 ;
  assign n28609 = n28607 & ~n28608 ;
  assign n28610 = n28550 ^ x300 ;
  assign n28611 = n28609 & ~n28610 ;
  assign n28612 = n28562 ^ x299 ;
  assign n28613 = ~n28611 & n28612 ;
  assign n28614 = n28574 ^ x298 ;
  assign n28615 = ~n28613 & n28614 ;
  assign n28988 = n28587 & ~n28615 ;
  assign n28989 = n28894 ^ x296 ;
  assign n28990 = n28988 & n28989 ;
  assign n28991 = n28896 ^ x311 ;
  assign n28992 = n28991 ^ n28897 ;
  assign n28993 = ~n28990 & n28992 ;
  assign n28994 = n28904 ^ x310 ;
  assign n28995 = n28993 & ~n28994 ;
  assign n28996 = n28910 ^ x309 ;
  assign n28997 = ~n28995 & n28996 ;
  assign n28998 = ~n28987 & ~n28997 ;
  assign n28999 = n28923 ^ x307 ;
  assign n29000 = ~n28998 & ~n28999 ;
  assign n29001 = n28930 ^ x306 ;
  assign n29002 = ~n29000 & n29001 ;
  assign n29003 = n28937 ^ x305 ;
  assign n29004 = ~n29002 & n29003 ;
  assign n29628 = n29005 ^ n29004 ;
  assign n28755 = n28247 ^ n28246 ;
  assign n28628 = n28243 ^ n28242 ;
  assign n28629 = n28628 ^ n28225 ;
  assign n28737 = n28736 ^ n28239 ;
  assign n28738 = n28631 & n28737 ;
  assign n28739 = n28738 ^ n28047 ;
  assign n28630 = n28241 ^ n28239 ;
  assign n28740 = n28739 ^ n28630 ;
  assign n28741 = n28628 ^ n28210 ;
  assign n28742 = n28741 ^ n28630 ;
  assign n28743 = n28742 ^ n28628 ;
  assign n28744 = n28740 & ~n28743 ;
  assign n28745 = n28744 ^ n28741 ;
  assign n28746 = n28629 & n28745 ;
  assign n28747 = n28746 ^ n28225 ;
  assign n28627 = n28245 ^ n28244 ;
  assign n28748 = n28747 ^ n28627 ;
  assign n28750 = n28409 ^ n28378 ;
  assign n28749 = n28747 ^ n28409 ;
  assign n28751 = n28750 ^ n28749 ;
  assign n28752 = n28748 & ~n28751 ;
  assign n28753 = n28752 ^ n28750 ;
  assign n28839 = n28755 ^ n28753 ;
  assign n29648 = n29628 ^ n28839 ;
  assign n29619 = n29003 ^ n29002 ;
  assign n29618 = n28748 ^ n28378 ;
  assign n29620 = n29619 ^ n29618 ;
  assign n29493 = n28997 ^ n28987 ;
  assign n29425 = n28996 ^ n28995 ;
  assign n29423 = n28712 ^ n27900 ;
  assign n29424 = n29423 ^ n28732 ;
  assign n29426 = n29425 ^ n29424 ;
  assign n29142 = n28424 ^ n28023 ;
  assign n29139 = n28398 ^ n28013 ;
  assign n29143 = n29142 ^ n29139 ;
  assign n29136 = n28614 ^ n28613 ;
  assign n29124 = n28291 ^ n28006 ;
  assign n29125 = n29124 ^ n28369 ;
  assign n29137 = n29136 ^ n29125 ;
  assign n28620 = n28363 ^ n27913 ;
  assign n28621 = n28620 ^ n28294 ;
  assign n28617 = n28608 ^ n28607 ;
  assign n28622 = n28621 ^ n28617 ;
  assign n28625 = n28606 ^ n28605 ;
  assign n29120 = n28625 ^ n28621 ;
  assign n28623 = n28360 ^ n27917 ;
  assign n28624 = n28623 ^ n28296 ;
  assign n28626 = n28625 ^ n28624 ;
  assign n29106 = n28357 ^ n27921 ;
  assign n29107 = n29106 ^ n28298 ;
  assign n29117 = n29107 ^ n28625 ;
  assign n29048 = n28333 ^ n27946 ;
  assign n29049 = n29048 ^ n28314 ;
  assign n29025 = n28330 ^ n27964 ;
  assign n29026 = n29025 ^ n28316 ;
  assign n28886 = n28885 ^ x304 ;
  assign n28943 = n28886 & ~n28942 ;
  assign n28944 = n28943 ^ x304 ;
  assign n28816 = n28815 ^ n28768 ;
  assign n28817 = n28630 ^ n28210 ;
  assign n28818 = n28817 ^ n28739 ;
  assign n28819 = n28818 ^ n28210 ;
  assign n28820 = n28819 ^ n27449 ;
  assign n28821 = n28820 ^ n26823 ;
  assign n28822 = n28821 ^ n28768 ;
  assign n28823 = n28822 ^ n28820 ;
  assign n28824 = ~n28816 & n28823 ;
  assign n28825 = n28824 ^ n28821 ;
  assign n28883 = n28825 ^ n26831 ;
  assign n28945 = n28944 ^ n28883 ;
  assign n28827 = n28224 ^ n26831 ;
  assign n28828 = n28827 ^ n28745 ;
  assign n28826 = n28820 ^ n28224 ;
  assign n28829 = n28828 ^ n28826 ;
  assign n28830 = n28829 ^ n28745 ;
  assign n28831 = n28825 & ~n28830 ;
  assign n28832 = n28831 ^ n28828 ;
  assign n28946 = n28832 ^ n26963 ;
  assign n28947 = n28946 ^ x319 ;
  assign n28948 = n28947 ^ n28883 ;
  assign n28949 = n28948 ^ n28946 ;
  assign n28950 = n28945 & ~n28949 ;
  assign n28951 = n28950 ^ n28947 ;
  assign n28765 = n28745 ^ n27309 ;
  assign n28833 = n28765 & n28832 ;
  assign n28763 = n28748 ^ n28371 ;
  assign n28764 = n28763 ^ n26963 ;
  assign n28834 = n28833 ^ n28764 ;
  assign n28952 = n28834 ^ n26983 ;
  assign n28954 = n28952 ^ x318 ;
  assign n28953 = n28952 ^ n28946 ;
  assign n28955 = n28954 ^ n28953 ;
  assign n28956 = ~n28951 & n28955 ;
  assign n28957 = n28956 ^ n28954 ;
  assign n28840 = n28839 ^ n28409 ;
  assign n28841 = n28840 ^ n27475 ;
  assign n28835 = n28748 ^ n27315 ;
  assign n28836 = ~n28834 & ~n28835 ;
  assign n28837 = n28836 ^ n26983 ;
  assign n28838 = n28837 ^ n27005 ;
  assign n28958 = n28841 ^ n28838 ;
  assign n28960 = n28958 ^ x317 ;
  assign n28959 = n28958 ^ n28952 ;
  assign n28961 = n28960 ^ n28959 ;
  assign n28962 = ~n28957 & n28961 ;
  assign n28963 = n28962 ^ n28960 ;
  assign n28842 = n28841 ^ n28837 ;
  assign n28843 = n28838 & ~n28842 ;
  assign n28844 = n28843 ^ n27005 ;
  assign n28964 = n28844 ^ n27024 ;
  assign n28754 = n28249 ^ n28248 ;
  assign n28757 = n28754 ^ n28409 ;
  assign n28756 = n28755 ^ n28754 ;
  assign n28758 = n28757 ^ n28756 ;
  assign n28759 = ~n28753 & n28758 ;
  assign n28760 = n28759 ^ n28757 ;
  assign n28761 = n28760 ^ n27488 ;
  assign n28965 = n28964 ^ n28761 ;
  assign n28967 = n28965 ^ x316 ;
  assign n28966 = n28965 ^ n28958 ;
  assign n28968 = n28967 ^ n28966 ;
  assign n28969 = ~n28963 & n28968 ;
  assign n28970 = n28969 ^ n28967 ;
  assign n28762 = n28761 ^ n27024 ;
  assign n28845 = n28844 ^ n28761 ;
  assign n28846 = n28762 & ~n28845 ;
  assign n28847 = n28846 ^ n27024 ;
  assign n28971 = n28847 ^ n27043 ;
  assign n28853 = n28251 ^ n28250 ;
  assign n28849 = n28662 ^ n28643 ;
  assign n28848 = n28754 ^ n28662 ;
  assign n28850 = n28849 ^ n28848 ;
  assign n28851 = n28760 & ~n28850 ;
  assign n28852 = n28851 ^ n28849 ;
  assign n28854 = n28853 ^ n28852 ;
  assign n28855 = n28854 ^ n28662 ;
  assign n28856 = n28855 ^ n27501 ;
  assign n28972 = n28971 ^ n28856 ;
  assign n28974 = n28972 ^ x315 ;
  assign n28973 = n28972 ^ n28965 ;
  assign n28975 = n28974 ^ n28973 ;
  assign n28976 = ~n28970 & n28975 ;
  assign n28977 = n28976 ^ n28974 ;
  assign n28857 = n28856 ^ n28847 ;
  assign n28858 = n28856 ^ n27043 ;
  assign n28859 = n28857 & n28858 ;
  assign n28860 = n28859 ^ n27043 ;
  assign n28978 = n28860 ^ n27114 ;
  assign n28861 = n28253 ^ n28252 ;
  assign n28863 = n28861 ^ n28662 ;
  assign n28862 = n28861 ^ n28853 ;
  assign n28864 = n28863 ^ n28862 ;
  assign n28865 = ~n28852 & ~n28864 ;
  assign n28866 = n28865 ^ n28863 ;
  assign n28867 = n28866 ^ n27514 ;
  assign n28979 = n28978 ^ n28867 ;
  assign n28981 = n28979 ^ x314 ;
  assign n28980 = n28979 ^ n28972 ;
  assign n28982 = n28981 ^ n28980 ;
  assign n28983 = ~n28977 & n28982 ;
  assign n28984 = n28983 ^ n28981 ;
  assign n28986 = n28970 ^ x315 ;
  assign n29006 = n29004 & ~n29005 ;
  assign n29007 = n28944 ^ x319 ;
  assign n29008 = n29007 ^ n28883 ;
  assign n29009 = n29006 & n29008 ;
  assign n29010 = n28951 ^ x318 ;
  assign n29011 = ~n29009 & n29010 ;
  assign n29012 = n28957 ^ x317 ;
  assign n29013 = n29011 & n29012 ;
  assign n29014 = n28963 ^ x316 ;
  assign n29015 = ~n29013 & ~n29014 ;
  assign n29016 = ~n28986 & n29015 ;
  assign n29017 = n28977 ^ x314 ;
  assign n29018 = ~n29016 & n29017 ;
  assign n29019 = n29018 ^ n28979 ;
  assign n29022 = n28984 & n29019 ;
  assign n28985 = n28984 ^ n28979 ;
  assign n29020 = n29019 ^ n28985 ;
  assign n29021 = x313 & n29020 ;
  assign n29023 = n29022 ^ n29021 ;
  assign n28875 = n28861 ^ n28681 ;
  assign n28876 = ~n28866 & n28875 ;
  assign n28872 = n28722 ^ n28254 ;
  assign n28873 = n28872 ^ n28255 ;
  assign n28874 = n28873 ^ n28861 ;
  assign n28877 = n28876 ^ n28874 ;
  assign n28878 = n28877 ^ n28722 ;
  assign n28879 = n28878 ^ n27526 ;
  assign n28880 = n28879 ^ n27180 ;
  assign n28871 = n27114 ^ x312 ;
  assign n28881 = n28880 ^ n28871 ;
  assign n28868 = n28867 ^ n28860 ;
  assign n28869 = n28867 ^ n27114 ;
  assign n28870 = ~n28868 & n28869 ;
  assign n28882 = n28881 ^ n28870 ;
  assign n29024 = n29023 ^ n28882 ;
  assign n29027 = n29026 ^ n29024 ;
  assign n29030 = n28327 ^ n27958 ;
  assign n29031 = n29030 ^ n28318 ;
  assign n29044 = n29031 ^ n29026 ;
  assign n29028 = n28984 ^ x313 ;
  assign n29029 = n29028 ^ n29018 ;
  assign n29032 = n29031 ^ n29029 ;
  assign n29036 = n28324 ^ n28323 ;
  assign n29033 = n29015 ^ n28986 ;
  assign n29034 = n28426 ^ n27949 ;
  assign n29035 = n29033 & n29034 ;
  assign n29037 = n29036 ^ n29035 ;
  assign n29038 = n29017 ^ n29016 ;
  assign n29039 = n29038 ^ n29035 ;
  assign n29040 = n29037 & n29039 ;
  assign n29041 = n29040 ^ n29036 ;
  assign n29042 = n29041 ^ n29029 ;
  assign n29043 = ~n29032 & ~n29042 ;
  assign n29045 = n29044 ^ n29043 ;
  assign n29046 = n29027 & n29045 ;
  assign n29047 = n29046 ^ n29026 ;
  assign n29050 = n29049 ^ n29047 ;
  assign n29051 = n28336 ^ n27943 ;
  assign n29052 = n29051 ^ n28312 ;
  assign n29053 = n29052 ^ n28588 ;
  assign n29054 = n29053 ^ n29052 ;
  assign n29055 = n29054 ^ n29047 ;
  assign n29056 = n29050 & n29055 ;
  assign n29057 = n29056 ^ n29053 ;
  assign n29059 = n28339 ^ n27940 ;
  assign n29060 = n29059 ^ n28310 ;
  assign n29062 = n29060 ^ n29052 ;
  assign n29058 = n28590 ^ n28588 ;
  assign n29061 = n29060 ^ n29058 ;
  assign n29063 = n29062 ^ n29061 ;
  assign n29064 = n29057 & n29063 ;
  assign n29065 = n29064 ^ n29062 ;
  assign n29067 = n28342 ^ n27937 ;
  assign n29068 = n29067 ^ n28308 ;
  assign n29070 = n29068 ^ n29060 ;
  assign n29066 = n28592 ^ n28591 ;
  assign n29069 = n29068 ^ n29066 ;
  assign n29071 = n29070 ^ n29069 ;
  assign n29072 = n29065 & n29071 ;
  assign n29073 = n29072 ^ n29070 ;
  assign n29075 = n28345 ^ n27934 ;
  assign n29076 = n29075 ^ n28306 ;
  assign n29078 = n29076 ^ n29068 ;
  assign n29074 = n28594 ^ n28593 ;
  assign n29077 = n29076 ^ n29074 ;
  assign n29079 = n29078 ^ n29077 ;
  assign n29080 = n29073 & n29079 ;
  assign n29081 = n29080 ^ n29078 ;
  assign n29083 = n28348 ^ n27931 ;
  assign n29084 = n29083 ^ n28304 ;
  assign n29086 = n29084 ^ n29076 ;
  assign n29082 = n28596 ^ n28595 ;
  assign n29085 = n29084 ^ n29082 ;
  assign n29087 = n29086 ^ n29085 ;
  assign n29088 = n29081 & ~n29087 ;
  assign n29089 = n29088 ^ n29086 ;
  assign n29091 = n28351 ^ n27928 ;
  assign n29092 = n29091 ^ n28302 ;
  assign n29094 = n29092 ^ n29084 ;
  assign n29090 = n28598 ^ n28597 ;
  assign n29093 = n29092 ^ n29090 ;
  assign n29095 = n29094 ^ n29093 ;
  assign n29096 = ~n29089 & ~n29095 ;
  assign n29097 = n29096 ^ n29094 ;
  assign n29099 = n28354 ^ n27925 ;
  assign n29100 = n29099 ^ n28300 ;
  assign n29102 = n29100 ^ n29092 ;
  assign n29098 = n28600 ^ n28599 ;
  assign n29101 = n29100 ^ n29098 ;
  assign n29103 = n29102 ^ n29101 ;
  assign n29104 = n29097 & ~n29103 ;
  assign n29105 = n29104 ^ n29102 ;
  assign n29110 = n29107 ^ n29100 ;
  assign n29108 = n28602 ^ n28601 ;
  assign n29109 = n29108 ^ n29107 ;
  assign n29111 = n29110 ^ n29109 ;
  assign n29112 = ~n29105 & ~n29111 ;
  assign n29113 = n29112 ^ n29110 ;
  assign n29114 = n28604 ^ n28603 ;
  assign n29115 = n29114 ^ n29107 ;
  assign n29116 = n29113 & ~n29115 ;
  assign n29118 = n29117 ^ n29116 ;
  assign n29119 = ~n28626 & n29118 ;
  assign n29121 = n29120 ^ n29119 ;
  assign n29122 = n28622 & ~n29121 ;
  assign n28618 = n28610 ^ n28609 ;
  assign n28619 = n28618 ^ n28617 ;
  assign n29123 = n29122 ^ n28619 ;
  assign n29127 = n28366 ^ n28002 ;
  assign n29128 = n29127 ^ n28292 ;
  assign n29129 = n29128 ^ n29125 ;
  assign n29126 = n29125 ^ n28618 ;
  assign n29130 = n29129 ^ n29126 ;
  assign n29131 = n29123 & n29130 ;
  assign n29132 = n29131 ^ n29126 ;
  assign n29133 = n28612 ^ n28611 ;
  assign n29134 = n29133 ^ n29125 ;
  assign n29135 = ~n29132 & n29134 ;
  assign n29138 = n29137 ^ n29135 ;
  assign n29140 = n29139 ^ n29136 ;
  assign n29141 = n29138 & ~n29140 ;
  assign n29144 = n29143 ^ n29141 ;
  assign n29261 = n28703 ^ n27909 ;
  assign n29262 = n29261 ^ n28699 ;
  assign n29263 = n29262 ^ n29142 ;
  assign n29264 = n29263 ^ n29262 ;
  assign n28616 = n28615 ^ n28587 ;
  assign n29265 = n29264 ^ n28616 ;
  assign n29266 = n29144 & n29265 ;
  assign n29267 = n29266 ^ n29263 ;
  assign n29274 = n28706 ^ n27906 ;
  assign n29275 = n29274 ^ n28697 ;
  assign n29277 = n29275 ^ n29262 ;
  assign n29268 = n28989 ^ n28988 ;
  assign n29276 = n29275 ^ n29268 ;
  assign n29278 = n29277 ^ n29276 ;
  assign n29279 = ~n29267 & n29278 ;
  assign n29280 = n29279 ^ n29277 ;
  assign n29285 = n28709 ^ n27903 ;
  assign n29286 = n29285 ^ n28695 ;
  assign n29288 = n29286 ^ n29275 ;
  assign n29281 = n28992 ^ n28990 ;
  assign n29287 = n29286 ^ n29281 ;
  assign n29289 = n29288 ^ n29287 ;
  assign n29290 = ~n29280 & ~n29289 ;
  assign n29291 = n29290 ^ n29288 ;
  assign n29292 = n28994 ^ n28993 ;
  assign n29427 = n29292 ^ n29286 ;
  assign n29428 = n29291 & ~n29427 ;
  assign n29429 = n29428 ^ n29286 ;
  assign n29490 = n29429 ^ n29425 ;
  assign n29491 = ~n29426 & n29490 ;
  assign n29492 = n29491 ^ n29429 ;
  assign n29521 = n29493 ^ n29492 ;
  assign n29522 = n28999 ^ n28998 ;
  assign n29523 = n29522 ^ n28766 ;
  assign n29524 = n29523 ^ n29522 ;
  assign n29525 = n29524 ^ n29492 ;
  assign n29526 = ~n29521 & n29525 ;
  assign n29527 = n29526 ^ n29523 ;
  assign n29569 = n29001 ^ n29000 ;
  assign n29571 = n29569 ^ n28818 ;
  assign n29570 = n29569 ^ n29522 ;
  assign n29572 = n29571 ^ n29570 ;
  assign n29573 = n29527 & ~n29572 ;
  assign n29574 = n29573 ^ n29571 ;
  assign n29575 = n28745 ^ n28225 ;
  assign n29622 = n29575 ^ n29569 ;
  assign n29623 = n29574 & n29622 ;
  assign n29621 = n29619 ^ n29575 ;
  assign n29624 = n29623 ^ n29621 ;
  assign n29625 = n29620 & ~n29624 ;
  assign n29626 = n29625 ^ n29619 ;
  assign n29649 = n29648 ^ n29626 ;
  assign n29650 = n29649 ^ n28840 ;
  assign n29638 = n29624 ^ n29618 ;
  assign n29639 = n29638 ^ n28748 ;
  assign n29640 = n29639 ^ n28371 ;
  assign n29576 = n29575 ^ n29574 ;
  assign n29577 = n29576 ^ n28745 ;
  assign n29578 = n29577 ^ n28224 ;
  assign n29494 = n29493 ^ n28766 ;
  assign n29495 = n29494 ^ n29492 ;
  assign n29496 = n29495 ^ n28767 ;
  assign n29430 = n29429 ^ n29426 ;
  assign n29431 = n29430 ^ n28733 ;
  assign n29432 = n29431 ^ n27319 ;
  assign n29282 = n29281 ^ n29280 ;
  assign n29283 = n29282 ^ n28707 ;
  assign n29145 = n29144 ^ n28616 ;
  assign n29146 = n29145 ^ n28424 ;
  assign n29147 = n29146 ^ n27250 ;
  assign n29236 = n29128 ^ n29123 ;
  assign n29237 = n29236 ^ n28367 ;
  assign n29148 = n29058 ^ n29057 ;
  assign n29149 = n29148 ^ n28337 ;
  assign n29150 = n29149 ^ n27806 ;
  assign n29172 = n29049 ^ n28588 ;
  assign n29173 = n29172 ^ n29047 ;
  assign n29174 = n29173 ^ n28334 ;
  assign n29151 = n29033 ^ n28320 ;
  assign n29152 = n27827 & ~n29151 ;
  assign n29153 = n29152 ^ n27825 ;
  assign n29154 = n29038 ^ n29037 ;
  assign n29155 = n29154 ^ n28325 ;
  assign n29156 = n29155 ^ n29152 ;
  assign n29157 = n29153 & ~n29156 ;
  assign n29158 = n29157 ^ n27825 ;
  assign n29159 = n29158 ^ n27820 ;
  assign n29160 = n29041 ^ n29031 ;
  assign n29161 = n29160 ^ n29029 ;
  assign n29162 = n29161 ^ n28328 ;
  assign n29163 = n29162 ^ n29158 ;
  assign n29164 = n29159 & ~n29163 ;
  assign n29165 = n29164 ^ n27820 ;
  assign n29166 = n29165 ^ n27815 ;
  assign n29167 = n29045 ^ n29024 ;
  assign n29168 = n29167 ^ n28331 ;
  assign n29169 = n29168 ^ n29165 ;
  assign n29170 = n29166 & n29169 ;
  assign n29171 = n29170 ^ n27815 ;
  assign n29175 = n29174 ^ n29171 ;
  assign n29176 = n29174 ^ n27810 ;
  assign n29177 = n29175 & n29176 ;
  assign n29178 = n29177 ^ n27810 ;
  assign n29179 = n29178 ^ n29149 ;
  assign n29180 = n29150 & n29179 ;
  assign n29181 = n29180 ^ n27806 ;
  assign n29182 = n29181 ^ n27802 ;
  assign n29183 = n29066 ^ n29065 ;
  assign n29184 = n29183 ^ n28340 ;
  assign n29185 = n29184 ^ n29181 ;
  assign n29186 = n29182 & n29185 ;
  assign n29187 = n29186 ^ n27802 ;
  assign n29188 = n29187 ^ n27798 ;
  assign n29189 = n29074 ^ n29073 ;
  assign n29190 = n29189 ^ n28343 ;
  assign n29191 = n29190 ^ n29187 ;
  assign n29192 = ~n29188 & n29191 ;
  assign n29193 = n29192 ^ n27798 ;
  assign n29194 = n29193 ^ n27794 ;
  assign n29195 = n29082 ^ n29081 ;
  assign n29196 = n29195 ^ n28346 ;
  assign n29197 = n29196 ^ n29193 ;
  assign n29198 = ~n29194 & ~n29197 ;
  assign n29199 = n29198 ^ n27794 ;
  assign n29200 = n29199 ^ n27789 ;
  assign n29201 = n29090 ^ n29089 ;
  assign n29202 = n29201 ^ n28349 ;
  assign n29203 = n29202 ^ n29199 ;
  assign n29204 = ~n29200 & n29203 ;
  assign n29205 = n29204 ^ n27789 ;
  assign n29206 = n29205 ^ n27787 ;
  assign n29207 = n29098 ^ n29097 ;
  assign n29208 = n29207 ^ n28352 ;
  assign n29209 = n29208 ^ n29205 ;
  assign n29210 = n29206 & n29209 ;
  assign n29211 = n29210 ^ n27787 ;
  assign n29212 = n29211 ^ n27347 ;
  assign n29213 = n29108 ^ n29105 ;
  assign n29214 = n29213 ^ n28355 ;
  assign n29215 = n29214 ^ n29211 ;
  assign n29216 = ~n29212 & ~n29215 ;
  assign n29217 = n29216 ^ n27347 ;
  assign n29218 = n29217 ^ n27344 ;
  assign n29219 = n29114 ^ n29113 ;
  assign n29220 = n29219 ^ n28358 ;
  assign n29221 = n29220 ^ n29217 ;
  assign n29222 = ~n29218 & n29221 ;
  assign n29223 = n29222 ^ n27344 ;
  assign n29224 = n29223 ^ n27340 ;
  assign n29225 = n29118 ^ n28624 ;
  assign n29226 = n29225 ^ n28361 ;
  assign n29227 = n29226 ^ n29223 ;
  assign n29228 = ~n29224 & ~n29227 ;
  assign n29229 = n29228 ^ n27340 ;
  assign n29230 = n29229 ^ n27336 ;
  assign n29231 = n29121 ^ n28617 ;
  assign n29232 = n29231 ^ n28364 ;
  assign n29233 = n29232 ^ n29229 ;
  assign n29234 = ~n29230 & ~n29233 ;
  assign n29235 = n29234 ^ n27336 ;
  assign n29238 = n29237 ^ n29235 ;
  assign n29239 = n29133 ^ n29132 ;
  assign n29240 = n29239 ^ n28370 ;
  assign n29241 = n29240 ^ n27408 ;
  assign n29242 = n29241 ^ n29235 ;
  assign n29243 = n29242 ^ n29240 ;
  assign n29244 = ~n29238 & n29243 ;
  assign n29245 = n29244 ^ n29241 ;
  assign n29246 = n29139 ^ n29138 ;
  assign n29247 = n29246 ^ n28398 ;
  assign n29249 = n29247 ^ n27279 ;
  assign n29248 = n29247 ^ n29240 ;
  assign n29250 = n29249 ^ n29248 ;
  assign n29251 = n29245 & n29250 ;
  assign n29252 = n29251 ^ n29249 ;
  assign n29254 = n29146 ^ n27876 ;
  assign n29253 = n29247 ^ n29146 ;
  assign n29255 = n29254 ^ n29253 ;
  assign n29256 = ~n29252 & n29255 ;
  assign n29257 = n29256 ^ n29254 ;
  assign n29258 = n29147 & ~n29257 ;
  assign n29259 = n29258 ^ n27250 ;
  assign n29260 = n29259 ^ n27241 ;
  assign n29269 = n29268 ^ n29267 ;
  assign n29270 = n29269 ^ n28704 ;
  assign n29271 = n29270 ^ n29259 ;
  assign n29272 = ~n29260 & n29271 ;
  assign n29273 = n29272 ^ n27241 ;
  assign n29284 = n29283 ^ n29273 ;
  assign n29293 = n29292 ^ n29291 ;
  assign n29294 = n29293 ^ n28710 ;
  assign n29295 = n29294 ^ n27248 ;
  assign n29296 = n29295 ^ n29273 ;
  assign n29297 = n29296 ^ n29294 ;
  assign n29298 = ~n29284 & n29297 ;
  assign n29299 = n29298 ^ n29295 ;
  assign n29420 = n29294 ^ n27323 ;
  assign n29421 = n29299 & ~n29420 ;
  assign n29422 = n29421 ^ n27323 ;
  assign n29486 = n29431 ^ n29422 ;
  assign n29487 = n29432 & n29486 ;
  assign n29488 = n29487 ^ n27319 ;
  assign n29520 = n29496 ^ n29488 ;
  assign n29528 = n29527 ^ n28818 ;
  assign n29529 = n29528 ^ n28819 ;
  assign n29530 = n29529 ^ n27444 ;
  assign n29531 = n29530 ^ n29488 ;
  assign n29532 = n29531 ^ n29529 ;
  assign n29533 = n29520 & ~n29532 ;
  assign n29534 = n29533 ^ n29530 ;
  assign n29566 = n29529 ^ n27449 ;
  assign n29567 = n29534 & n29566 ;
  assign n29568 = n29567 ^ n27449 ;
  assign n29641 = n29577 ^ n29568 ;
  assign n29642 = ~n29578 & n29641 ;
  assign n29643 = n29642 ^ n28224 ;
  assign n29644 = n29643 ^ n29639 ;
  assign n29645 = n29640 & ~n29644 ;
  assign n29646 = n29645 ^ n28371 ;
  assign n29647 = n29646 ^ n27475 ;
  assign n29656 = n29650 ^ n29647 ;
  assign n29692 = n29656 ^ x412 ;
  assign n29657 = n29643 ^ n29640 ;
  assign n29658 = n29657 ^ x413 ;
  assign n29579 = n29578 ^ n29568 ;
  assign n29535 = n29534 ^ n27449 ;
  assign n29536 = n29535 ^ x415 ;
  assign n29301 = n29273 ^ n27248 ;
  assign n29302 = n29301 ^ n29283 ;
  assign n29303 = n29302 ^ x403 ;
  assign n29304 = n29257 ^ n27250 ;
  assign n29305 = n29304 ^ x405 ;
  assign n29396 = n29245 ^ n27279 ;
  assign n29306 = n29235 ^ n27408 ;
  assign n29307 = n29306 ^ n29237 ;
  assign n29308 = n29307 ^ x392 ;
  assign n29310 = n29171 ^ n27810 ;
  assign n29311 = n29310 ^ n29174 ;
  assign n29312 = n29311 ^ x387 ;
  assign n29314 = n29033 ^ n27828 ;
  assign n29315 = x391 & ~n29314 ;
  assign n29316 = n29315 ^ x390 ;
  assign n29317 = n29156 ^ n27825 ;
  assign n29318 = n29317 ^ n29315 ;
  assign n29319 = n29316 & ~n29318 ;
  assign n29320 = n29319 ^ x390 ;
  assign n29321 = n29320 ^ x389 ;
  assign n29322 = n29162 ^ n29159 ;
  assign n29323 = n29322 ^ n29320 ;
  assign n29324 = n29321 & ~n29323 ;
  assign n29325 = n29324 ^ x389 ;
  assign n29313 = n29168 ^ n29166 ;
  assign n29326 = n29325 ^ n29313 ;
  assign n29328 = n29311 ^ x388 ;
  assign n29327 = n29325 ^ n29311 ;
  assign n29329 = n29328 ^ n29327 ;
  assign n29330 = n29326 & n29329 ;
  assign n29331 = n29330 ^ n29328 ;
  assign n29332 = n29312 & ~n29331 ;
  assign n29333 = n29332 ^ x387 ;
  assign n29334 = n29333 ^ x386 ;
  assign n29335 = n29178 ^ n27806 ;
  assign n29336 = n29335 ^ n29149 ;
  assign n29337 = n29336 ^ n29333 ;
  assign n29338 = n29334 & n29337 ;
  assign n29339 = n29338 ^ x386 ;
  assign n29309 = n29184 ^ n29182 ;
  assign n29340 = n29339 ^ n29309 ;
  assign n29341 = n29190 ^ n29188 ;
  assign n29342 = n29341 ^ x385 ;
  assign n29343 = n29342 ^ n29339 ;
  assign n29344 = n29343 ^ n29341 ;
  assign n29345 = n29340 & n29344 ;
  assign n29346 = n29345 ^ n29342 ;
  assign n29347 = n29196 ^ n29194 ;
  assign n29349 = n29347 ^ x384 ;
  assign n29348 = n29347 ^ n29341 ;
  assign n29350 = n29349 ^ n29348 ;
  assign n29351 = ~n29346 & n29350 ;
  assign n29352 = n29351 ^ n29349 ;
  assign n29353 = n29202 ^ n29200 ;
  assign n29355 = n29353 ^ x399 ;
  assign n29354 = n29353 ^ n29347 ;
  assign n29356 = n29355 ^ n29354 ;
  assign n29357 = ~n29352 & n29356 ;
  assign n29358 = n29357 ^ n29355 ;
  assign n29359 = n29208 ^ n29206 ;
  assign n29361 = n29359 ^ x398 ;
  assign n29360 = n29359 ^ n29353 ;
  assign n29362 = n29361 ^ n29360 ;
  assign n29363 = ~n29358 & n29362 ;
  assign n29364 = n29363 ^ n29361 ;
  assign n29365 = n29214 ^ n29212 ;
  assign n29367 = n29365 ^ x397 ;
  assign n29366 = n29365 ^ n29359 ;
  assign n29368 = n29367 ^ n29366 ;
  assign n29369 = ~n29364 & n29368 ;
  assign n29370 = n29369 ^ n29367 ;
  assign n29371 = n29220 ^ n29218 ;
  assign n29373 = n29371 ^ x396 ;
  assign n29372 = n29371 ^ n29365 ;
  assign n29374 = n29373 ^ n29372 ;
  assign n29375 = ~n29370 & n29374 ;
  assign n29376 = n29375 ^ n29373 ;
  assign n29377 = n29226 ^ n29224 ;
  assign n29379 = n29377 ^ x395 ;
  assign n29378 = n29377 ^ n29371 ;
  assign n29380 = n29379 ^ n29378 ;
  assign n29381 = ~n29376 & n29380 ;
  assign n29382 = n29381 ^ n29379 ;
  assign n29383 = n29232 ^ n29230 ;
  assign n29385 = n29383 ^ x394 ;
  assign n29384 = n29383 ^ n29377 ;
  assign n29386 = n29385 ^ n29384 ;
  assign n29387 = ~n29382 & n29386 ;
  assign n29388 = n29387 ^ n29385 ;
  assign n29390 = n29307 ^ x393 ;
  assign n29389 = n29383 ^ n29307 ;
  assign n29391 = n29390 ^ n29389 ;
  assign n29392 = n29388 & ~n29391 ;
  assign n29393 = n29392 ^ n29390 ;
  assign n29394 = ~n29308 & n29393 ;
  assign n29395 = n29394 ^ x392 ;
  assign n29397 = n29396 ^ n29395 ;
  assign n29398 = n29252 ^ n27876 ;
  assign n29399 = n29398 ^ x407 ;
  assign n29400 = n29399 ^ n29395 ;
  assign n29401 = n29400 ^ n29398 ;
  assign n29402 = n29397 & n29401 ;
  assign n29403 = n29402 ^ n29399 ;
  assign n29405 = n29304 ^ x406 ;
  assign n29404 = n29398 ^ n29304 ;
  assign n29406 = n29405 ^ n29404 ;
  assign n29407 = ~n29403 & n29406 ;
  assign n29408 = n29407 ^ n29405 ;
  assign n29409 = n29305 & ~n29408 ;
  assign n29410 = n29409 ^ x405 ;
  assign n29411 = n29410 ^ x404 ;
  assign n29412 = n29270 ^ n29260 ;
  assign n29413 = n29412 ^ n29410 ;
  assign n29414 = n29411 & ~n29413 ;
  assign n29415 = n29414 ^ x404 ;
  assign n29416 = n29415 ^ n29302 ;
  assign n29417 = ~n29303 & n29416 ;
  assign n29418 = n29417 ^ x403 ;
  assign n29300 = n29299 ^ n27323 ;
  assign n29419 = n29418 ^ n29300 ;
  assign n29433 = n29432 ^ n29422 ;
  assign n29434 = n29433 ^ x402 ;
  assign n29435 = n29434 ^ n29300 ;
  assign n29436 = n29435 ^ n29433 ;
  assign n29437 = ~n29419 & n29436 ;
  assign n29438 = n29437 ^ n29434 ;
  assign n29489 = n29488 ^ n27444 ;
  assign n29497 = n29496 ^ n29489 ;
  assign n29499 = n29497 ^ x401 ;
  assign n29498 = n29497 ^ n29433 ;
  assign n29500 = n29499 ^ n29498 ;
  assign n29501 = n29438 & ~n29500 ;
  assign n29502 = n29501 ^ n29499 ;
  assign n29517 = n29497 ^ x400 ;
  assign n29518 = ~n29502 & n29517 ;
  assign n29519 = n29518 ^ x400 ;
  assign n29562 = n29535 ^ n29519 ;
  assign n29563 = ~n29536 & n29562 ;
  assign n29564 = n29563 ^ x415 ;
  assign n29659 = n29579 ^ n29564 ;
  assign n29660 = n29657 ^ x414 ;
  assign n29661 = n29660 ^ n29657 ;
  assign n29662 = n29661 ^ n29564 ;
  assign n29663 = n29659 & n29662 ;
  assign n29664 = n29663 ^ n29660 ;
  assign n29665 = n29658 & ~n29664 ;
  assign n29666 = n29665 ^ x413 ;
  assign n29693 = n29692 ^ n29666 ;
  assign n29565 = n29564 ^ x414 ;
  assign n29580 = n29579 ^ n29565 ;
  assign n29537 = n29536 ^ n29519 ;
  assign n29439 = n29438 ^ x401 ;
  assign n29440 = n29300 ^ x402 ;
  assign n29441 = n29440 ^ n29418 ;
  assign n29442 = n29382 ^ x394 ;
  assign n29443 = n29314 ^ x391 ;
  assign n29444 = n29318 ^ x390 ;
  assign n29445 = ~n29443 & n29444 ;
  assign n29446 = n29323 ^ x389 ;
  assign n29447 = ~n29445 & ~n29446 ;
  assign n29448 = n29326 ^ x388 ;
  assign n29449 = ~n29447 & ~n29448 ;
  assign n29450 = n29331 ^ x387 ;
  assign n29451 = n29449 & n29450 ;
  assign n29452 = n29337 ^ x386 ;
  assign n29453 = ~n29451 & n29452 ;
  assign n29454 = n29340 ^ x385 ;
  assign n29455 = n29453 & n29454 ;
  assign n29456 = n29346 ^ x384 ;
  assign n29457 = n29455 & ~n29456 ;
  assign n29458 = n29352 ^ x399 ;
  assign n29459 = n29457 & ~n29458 ;
  assign n29460 = n29358 ^ x398 ;
  assign n29461 = ~n29459 & n29460 ;
  assign n29462 = n29364 ^ x397 ;
  assign n29463 = n29461 & n29462 ;
  assign n29464 = n29370 ^ x396 ;
  assign n29465 = ~n29463 & ~n29464 ;
  assign n29466 = n29376 ^ x395 ;
  assign n29467 = n29465 & ~n29466 ;
  assign n29468 = n29442 & ~n29467 ;
  assign n29469 = n29388 ^ x393 ;
  assign n29470 = n29468 & ~n29469 ;
  assign n29471 = n29393 ^ x392 ;
  assign n29472 = ~n29470 & n29471 ;
  assign n29473 = n29395 ^ x407 ;
  assign n29474 = n29473 ^ n29396 ;
  assign n29475 = n29472 & n29474 ;
  assign n29476 = n29403 ^ x406 ;
  assign n29477 = n29475 & ~n29476 ;
  assign n29478 = n29408 ^ x405 ;
  assign n29479 = ~n29477 & n29478 ;
  assign n29480 = n29412 ^ n29411 ;
  assign n29481 = ~n29479 & ~n29480 ;
  assign n29482 = n29415 ^ n29303 ;
  assign n29483 = n29481 & n29482 ;
  assign n29484 = n29441 & ~n29483 ;
  assign n29485 = n29439 & ~n29484 ;
  assign n29503 = n29502 ^ x400 ;
  assign n29538 = n29485 & ~n29503 ;
  assign n29581 = ~n29537 & ~n29538 ;
  assign n29689 = n29580 & ~n29581 ;
  assign n29690 = n29664 ^ x413 ;
  assign n29691 = n29689 & ~n29690 ;
  assign n29723 = n29693 ^ n29691 ;
  assign n29724 = n29723 ^ n29183 ;
  assign n29725 = n29690 ^ n29689 ;
  assign n29726 = n29725 ^ n29148 ;
  assign n29582 = n29581 ^ n29580 ;
  assign n29539 = n29538 ^ n29537 ;
  assign n29505 = n29034 ^ n29033 ;
  assign n29506 = n29483 ^ n29441 ;
  assign n29507 = n29505 & ~n29506 ;
  assign n29508 = n29507 ^ n29154 ;
  assign n29509 = n29484 ^ n29439 ;
  assign n29510 = n29509 ^ n29507 ;
  assign n29511 = ~n29508 & ~n29510 ;
  assign n29512 = n29511 ^ n29154 ;
  assign n29504 = n29503 ^ n29485 ;
  assign n29513 = n29512 ^ n29504 ;
  assign n29514 = n29512 ^ n29161 ;
  assign n29515 = n29513 & n29514 ;
  assign n29516 = n29515 ^ n29161 ;
  assign n29540 = n29539 ^ n29516 ;
  assign n29559 = n29539 ^ n29167 ;
  assign n29560 = n29540 & ~n29559 ;
  assign n29561 = n29560 ^ n29167 ;
  assign n29583 = n29582 ^ n29561 ;
  assign n29727 = n29582 ^ n29173 ;
  assign n29728 = n29583 & n29727 ;
  assign n29729 = n29728 ^ n29173 ;
  assign n29730 = n29729 ^ n29725 ;
  assign n29731 = ~n29726 & ~n29730 ;
  assign n29732 = n29731 ^ n29148 ;
  assign n29733 = n29732 ^ n29723 ;
  assign n29734 = ~n29724 & n29733 ;
  assign n29735 = n29734 ^ n29183 ;
  assign n30291 = n29735 ^ n29189 ;
  assign n29667 = n29666 ^ n29656 ;
  assign n29651 = n29650 ^ n29646 ;
  assign n29652 = ~n29647 & ~n29651 ;
  assign n29653 = n29652 ^ n27475 ;
  assign n29633 = n29008 ^ n29006 ;
  assign n29632 = n28760 ^ n28643 ;
  assign n29634 = n29633 ^ n29632 ;
  assign n29627 = n29626 ^ n28839 ;
  assign n29629 = n29628 ^ n29626 ;
  assign n29630 = ~n29627 & ~n29629 ;
  assign n29631 = n29630 ^ n28839 ;
  assign n29635 = n29634 ^ n29631 ;
  assign n29636 = n29635 ^ n28760 ;
  assign n29637 = n29636 ^ n27488 ;
  assign n29654 = n29653 ^ n29637 ;
  assign n29668 = n29654 ^ x412 ;
  assign n29669 = n29668 ^ n29654 ;
  assign n29670 = n29669 ^ n29656 ;
  assign n29671 = n29667 & ~n29670 ;
  assign n29672 = n29671 ^ n29668 ;
  assign n29695 = n29672 ^ x411 ;
  assign n29694 = ~n29691 & ~n29693 ;
  assign n29721 = n29695 ^ n29694 ;
  assign n30292 = n30291 ^ n29721 ;
  assign n29784 = n29448 ^ n29447 ;
  assign n29899 = n29784 ^ n29231 ;
  assign n29616 = n29444 ^ n29443 ;
  assign n29617 = n29616 ^ n29219 ;
  assign n29696 = n29694 & n29695 ;
  assign n29684 = n29010 ^ n29009 ;
  assign n29682 = n29633 ^ n28854 ;
  assign n29680 = n29632 ^ n29631 ;
  assign n29681 = n29634 & ~n29680 ;
  assign n29683 = n29682 ^ n29681 ;
  assign n29685 = n29684 ^ n29683 ;
  assign n29686 = n29685 ^ n28855 ;
  assign n29676 = n29653 ^ n29636 ;
  assign n29677 = ~n29637 & n29676 ;
  assign n29678 = n29677 ^ n27488 ;
  assign n29679 = n29678 ^ n27501 ;
  assign n29687 = n29686 ^ n29679 ;
  assign n29655 = n29654 ^ x411 ;
  assign n29673 = n29655 & ~n29672 ;
  assign n29674 = n29673 ^ x411 ;
  assign n29675 = n29674 ^ x410 ;
  assign n29688 = n29687 ^ n29675 ;
  assign n29719 = n29696 ^ n29688 ;
  assign n29720 = n29719 ^ n29195 ;
  assign n29722 = n29721 ^ n29189 ;
  assign n29736 = n29735 ^ n29721 ;
  assign n29737 = ~n29722 & n29736 ;
  assign n29738 = n29737 ^ n29189 ;
  assign n29739 = n29738 ^ n29719 ;
  assign n29740 = n29720 & n29739 ;
  assign n29741 = n29740 ^ n29195 ;
  assign n29712 = n29687 ^ n29674 ;
  assign n29713 = n29687 ^ x410 ;
  assign n29714 = n29712 & ~n29713 ;
  assign n29715 = n29714 ^ x410 ;
  assign n29716 = n29715 ^ x409 ;
  assign n29706 = n29684 ^ n28854 ;
  assign n29707 = n29683 & n29706 ;
  assign n29708 = n29707 ^ n28854 ;
  assign n29704 = n29012 ^ n29011 ;
  assign n29703 = n28866 ^ n28681 ;
  assign n29705 = n29704 ^ n29703 ;
  assign n29709 = n29708 ^ n29705 ;
  assign n29710 = n29709 ^ n28866 ;
  assign n29698 = n29686 ^ n27501 ;
  assign n29699 = n29686 ^ n29678 ;
  assign n29700 = n29698 & ~n29699 ;
  assign n29701 = n29700 ^ n27501 ;
  assign n29702 = n29701 ^ n27514 ;
  assign n29711 = n29710 ^ n29702 ;
  assign n29717 = n29716 ^ n29711 ;
  assign n29697 = n29688 & ~n29696 ;
  assign n29718 = n29717 ^ n29697 ;
  assign n29742 = n29741 ^ n29718 ;
  assign n29756 = n29711 ^ n29697 ;
  assign n29759 = n29756 ^ n29715 ;
  assign n29760 = x409 & n29759 ;
  assign n29757 = n29715 ^ n29697 ;
  assign n29758 = n29756 & n29757 ;
  assign n29761 = n29760 ^ n29758 ;
  assign n29749 = n29708 ^ n29704 ;
  assign n29750 = ~n29705 & ~n29749 ;
  assign n29746 = n29013 ^ n28877 ;
  assign n29747 = n29746 ^ n29014 ;
  assign n29748 = n29747 ^ n29704 ;
  assign n29751 = n29750 ^ n29748 ;
  assign n29752 = n29751 ^ n28879 ;
  assign n29753 = n29752 ^ x408 ;
  assign n29754 = n29753 ^ n27514 ;
  assign n29743 = n29710 ^ n29701 ;
  assign n29744 = n29710 ^ n27514 ;
  assign n29745 = ~n29743 & ~n29744 ;
  assign n29755 = n29754 ^ n29745 ;
  assign n29762 = n29761 ^ n29755 ;
  assign n29763 = n29762 ^ n29201 ;
  assign n29764 = n29763 ^ n29718 ;
  assign n29765 = n29764 ^ n29762 ;
  assign n29766 = ~n29742 & n29765 ;
  assign n29767 = n29766 ^ n29763 ;
  assign n29769 = n29443 ^ n29207 ;
  assign n29768 = n29762 ^ n29443 ;
  assign n29770 = n29769 ^ n29768 ;
  assign n29771 = ~n29767 & ~n29770 ;
  assign n29772 = n29771 ^ n29769 ;
  assign n29774 = n29219 ^ n29213 ;
  assign n29773 = n29443 ^ n29219 ;
  assign n29775 = n29774 ^ n29773 ;
  assign n29776 = n29772 & ~n29775 ;
  assign n29777 = n29776 ^ n29774 ;
  assign n29778 = ~n29617 & ~n29777 ;
  assign n29779 = n29778 ^ n29219 ;
  assign n29615 = n29446 ^ n29445 ;
  assign n29780 = n29779 ^ n29615 ;
  assign n29781 = n29779 ^ n29225 ;
  assign n29782 = n29780 & n29781 ;
  assign n29783 = n29782 ^ n29225 ;
  assign n29900 = n29899 ^ n29783 ;
  assign n29901 = n29900 ^ n29231 ;
  assign n29902 = n29901 ^ n28621 ;
  assign n30124 = n29902 ^ n27913 ;
  assign n29903 = n29615 ^ n29225 ;
  assign n29904 = n29903 ^ n29779 ;
  assign n29905 = n29904 ^ n29225 ;
  assign n29906 = n29905 ^ n28624 ;
  assign n29907 = n29906 ^ n27917 ;
  assign n29908 = n29772 ^ n29100 ;
  assign n29909 = n29908 ^ n27925 ;
  assign n29910 = n29767 ^ n29092 ;
  assign n29911 = n29910 ^ n27928 ;
  assign n29912 = n29742 ^ n29084 ;
  assign n29913 = n29912 ^ n27931 ;
  assign n29914 = n29739 ^ n29076 ;
  assign n29915 = n29914 ^ n27934 ;
  assign n29584 = n29583 ^ n29049 ;
  assign n29917 = n29584 ^ n27946 ;
  assign n29541 = n29540 ^ n29026 ;
  assign n29542 = n29541 ^ n27964 ;
  assign n29543 = n29513 ^ n29031 ;
  assign n29544 = n29543 ^ n27958 ;
  assign n29545 = n29506 ^ n29034 ;
  assign n29546 = ~n28320 & ~n29545 ;
  assign n29547 = n29546 ^ n27952 ;
  assign n29548 = n29510 ^ n29036 ;
  assign n29549 = n29548 ^ n29546 ;
  assign n29550 = ~n29547 & ~n29549 ;
  assign n29551 = n29550 ^ n27952 ;
  assign n29552 = n29551 ^ n29543 ;
  assign n29553 = n29544 & n29552 ;
  assign n29554 = n29553 ^ n27958 ;
  assign n29555 = n29554 ^ n29541 ;
  assign n29556 = ~n29542 & ~n29555 ;
  assign n29557 = n29556 ^ n27964 ;
  assign n29918 = n29584 ^ n29557 ;
  assign n29919 = n29917 & ~n29918 ;
  assign n29920 = n29919 ^ n27946 ;
  assign n29921 = n29920 ^ n27943 ;
  assign n29922 = n29730 ^ n29052 ;
  assign n29923 = n29922 ^ n29920 ;
  assign n29924 = ~n29921 & ~n29923 ;
  assign n29925 = n29924 ^ n27943 ;
  assign n29916 = n29733 ^ n29060 ;
  assign n29926 = n29925 ^ n29916 ;
  assign n29927 = n29736 ^ n29068 ;
  assign n29928 = n29927 ^ n27940 ;
  assign n29929 = n29928 ^ n29916 ;
  assign n29930 = n29929 ^ n29927 ;
  assign n29931 = ~n29926 & ~n29930 ;
  assign n29932 = n29931 ^ n29928 ;
  assign n29934 = n29914 ^ n27937 ;
  assign n29933 = n29927 ^ n29914 ;
  assign n29935 = n29934 ^ n29933 ;
  assign n29936 = n29932 & ~n29935 ;
  assign n29937 = n29936 ^ n29934 ;
  assign n29938 = n29915 & n29937 ;
  assign n29939 = n29938 ^ n27934 ;
  assign n29940 = n29939 ^ n29912 ;
  assign n29941 = ~n29913 & ~n29940 ;
  assign n29942 = n29941 ^ n27931 ;
  assign n29943 = n29942 ^ n29910 ;
  assign n29944 = ~n29911 & n29943 ;
  assign n29945 = n29944 ^ n27928 ;
  assign n29946 = n29945 ^ n29908 ;
  assign n29947 = ~n29909 & n29946 ;
  assign n29948 = n29947 ^ n27925 ;
  assign n29949 = n29948 ^ n27921 ;
  assign n29950 = n29777 ^ n29616 ;
  assign n29951 = n29950 ^ n29219 ;
  assign n29952 = n29951 ^ n29107 ;
  assign n29953 = n29952 ^ n29948 ;
  assign n29954 = ~n29949 & ~n29953 ;
  assign n29955 = n29954 ^ n27921 ;
  assign n29956 = n29955 ^ n29906 ;
  assign n29957 = n29907 & n29956 ;
  assign n29958 = n29957 ^ n27917 ;
  assign n30125 = n30124 ^ n29958 ;
  assign n30069 = n29945 ^ n27925 ;
  assign n30070 = n30069 ^ n29908 ;
  assign n30071 = n30070 ^ x492 ;
  assign n30103 = n29942 ^ n27928 ;
  assign n30104 = n30103 ^ n29910 ;
  assign n30072 = n29939 ^ n27931 ;
  assign n30073 = n30072 ^ n29912 ;
  assign n30074 = n30073 ^ x494 ;
  assign n30075 = n29937 ^ n27934 ;
  assign n30076 = n30075 ^ x495 ;
  assign n30078 = n29916 ^ n27940 ;
  assign n30079 = n30078 ^ n29925 ;
  assign n30080 = n30079 ^ x481 ;
  assign n29586 = n29554 ^ n29542 ;
  assign n29587 = n29586 ^ x484 ;
  assign n29589 = n29506 ^ n28321 ;
  assign n29590 = x487 & n29589 ;
  assign n29591 = n29590 ^ x486 ;
  assign n29592 = n29548 ^ n29547 ;
  assign n29593 = n29592 ^ n29590 ;
  assign n29594 = n29591 & n29593 ;
  assign n29595 = n29594 ^ x486 ;
  assign n29588 = n29551 ^ n29544 ;
  assign n29596 = n29595 ^ n29588 ;
  assign n29597 = n29586 ^ x485 ;
  assign n29598 = n29597 ^ n29586 ;
  assign n29599 = n29598 ^ n29588 ;
  assign n29600 = n29596 & ~n29599 ;
  assign n29601 = n29600 ^ n29597 ;
  assign n29602 = ~n29587 & n29601 ;
  assign n29603 = n29602 ^ x484 ;
  assign n29604 = n29603 ^ x483 ;
  assign n29558 = n29557 ^ n27946 ;
  assign n29585 = n29584 ^ n29558 ;
  assign n30082 = n29603 ^ n29585 ;
  assign n30083 = n29604 & n30082 ;
  assign n30084 = n30083 ^ x483 ;
  assign n30081 = n29922 ^ n29921 ;
  assign n30085 = n30084 ^ n30081 ;
  assign n30086 = n30079 ^ x482 ;
  assign n30087 = n30086 ^ n30079 ;
  assign n30088 = n30087 ^ n30081 ;
  assign n30089 = ~n30085 & n30088 ;
  assign n30090 = n30089 ^ n30086 ;
  assign n30091 = ~n30080 & n30090 ;
  assign n30092 = n30091 ^ x481 ;
  assign n30077 = n29932 ^ n27937 ;
  assign n30093 = n30092 ^ n30077 ;
  assign n30094 = n30092 ^ x480 ;
  assign n30095 = ~n30093 & n30094 ;
  assign n30096 = n30095 ^ x480 ;
  assign n30097 = n30096 ^ n30075 ;
  assign n30098 = ~n30076 & n30097 ;
  assign n30099 = n30098 ^ x495 ;
  assign n30100 = n30099 ^ n30073 ;
  assign n30101 = ~n30074 & n30100 ;
  assign n30102 = n30101 ^ x494 ;
  assign n30105 = n30104 ^ n30102 ;
  assign n30106 = n30070 ^ x493 ;
  assign n30107 = n30106 ^ n30070 ;
  assign n30108 = n30107 ^ n30102 ;
  assign n30109 = ~n30105 & n30108 ;
  assign n30110 = n30109 ^ n30106 ;
  assign n30111 = n30071 & ~n30110 ;
  assign n30112 = n30111 ^ x492 ;
  assign n30113 = n30112 ^ x491 ;
  assign n30114 = n29952 ^ n29949 ;
  assign n30115 = n30114 ^ n30112 ;
  assign n30116 = n30113 & ~n30115 ;
  assign n30117 = n30116 ^ x491 ;
  assign n30118 = n30117 ^ x490 ;
  assign n30119 = n29955 ^ n27917 ;
  assign n30120 = n30119 ^ n29906 ;
  assign n30121 = n30120 ^ n30117 ;
  assign n30122 = n30118 & ~n30121 ;
  assign n30123 = n30122 ^ x490 ;
  assign n30126 = n30125 ^ n30123 ;
  assign n29959 = n29958 ^ n29902 ;
  assign n29960 = n29958 ^ n27913 ;
  assign n29961 = ~n29959 & ~n29960 ;
  assign n29962 = n29961 ^ n27913 ;
  assign n29785 = n29784 ^ n29783 ;
  assign n29613 = n29450 ^ n29449 ;
  assign n29786 = n29613 ^ n29231 ;
  assign n29787 = n29786 ^ n29613 ;
  assign n29788 = n29787 ^ n29783 ;
  assign n29789 = ~n29785 & ~n29788 ;
  assign n29790 = n29789 ^ n29786 ;
  assign n29897 = n29790 ^ n29128 ;
  assign n29898 = n29897 ^ n28002 ;
  assign n30127 = n29962 ^ n29898 ;
  assign n30128 = n30127 ^ x489 ;
  assign n30129 = n30128 ^ n30123 ;
  assign n30130 = n30129 ^ n30127 ;
  assign n30131 = ~n30126 & n30130 ;
  assign n30132 = n30131 ^ n30128 ;
  assign n29612 = n29452 ^ n29451 ;
  assign n29966 = n29612 ^ n29239 ;
  assign n29614 = n29613 ^ n29236 ;
  assign n29791 = ~n29614 & n29790 ;
  assign n29792 = n29791 ^ n29236 ;
  assign n29967 = n29966 ^ n29792 ;
  assign n29968 = n29967 ^ n29239 ;
  assign n29969 = n29968 ^ n29125 ;
  assign n30066 = n29969 ^ n28006 ;
  assign n29963 = n29962 ^ n29897 ;
  assign n29964 = ~n29898 & ~n29963 ;
  assign n29965 = n29964 ^ n28002 ;
  assign n30067 = n30066 ^ n29965 ;
  assign n30134 = n30067 ^ x488 ;
  assign n30133 = n30127 ^ n30067 ;
  assign n30135 = n30134 ^ n30133 ;
  assign n30136 = n30132 & ~n30135 ;
  assign n30137 = n30136 ^ n30134 ;
  assign n30219 = n30137 ^ x503 ;
  assign n30220 = n30090 ^ x481 ;
  assign n29605 = n29604 ^ n29585 ;
  assign n29606 = n29601 ^ x484 ;
  assign n30221 = n29605 & n29606 ;
  assign n30222 = n30081 ^ x482 ;
  assign n30223 = n30222 ^ n30084 ;
  assign n30224 = n30221 & ~n30223 ;
  assign n30225 = n30220 & n30224 ;
  assign n30226 = n30077 ^ x480 ;
  assign n30227 = n30226 ^ n30092 ;
  assign n30228 = n30225 & ~n30227 ;
  assign n30229 = n30096 ^ n30076 ;
  assign n30230 = ~n30228 & ~n30229 ;
  assign n30231 = n30099 ^ n30074 ;
  assign n30232 = n30230 & ~n30231 ;
  assign n30233 = n30104 ^ x493 ;
  assign n30234 = n30233 ^ n30102 ;
  assign n30235 = ~n30232 & ~n30234 ;
  assign n30236 = n30110 ^ x492 ;
  assign n30237 = n30235 & ~n30236 ;
  assign n30238 = n30114 ^ n30113 ;
  assign n30239 = n30237 & ~n30238 ;
  assign n30240 = n30120 ^ n30118 ;
  assign n30241 = n30239 & ~n30240 ;
  assign n30242 = n30125 ^ x489 ;
  assign n30243 = n30242 ^ n30123 ;
  assign n30244 = n30241 & ~n30243 ;
  assign n30245 = n30132 ^ x488 ;
  assign n30246 = ~n30244 & ~n30245 ;
  assign n30247 = ~n30219 & n30246 ;
  assign n30068 = n30067 ^ x503 ;
  assign n30138 = ~n30068 & n30137 ;
  assign n30139 = n30138 ^ x503 ;
  assign n29970 = n29969 ^ n29965 ;
  assign n29971 = n29138 ^ n28006 ;
  assign n29793 = n29792 ^ n29612 ;
  assign n29794 = n29246 ^ n29239 ;
  assign n29795 = n29794 ^ n29246 ;
  assign n29796 = n29795 ^ n29612 ;
  assign n29797 = n29793 & ~n29796 ;
  assign n29798 = n29797 ^ n29794 ;
  assign n29610 = n29454 ^ n29453 ;
  assign n29811 = n29798 ^ n29610 ;
  assign n29972 = n29971 ^ n29811 ;
  assign n29973 = n29972 ^ n29138 ;
  assign n29974 = n29973 ^ n29965 ;
  assign n29975 = n29974 ^ n29811 ;
  assign n29976 = ~n29970 & n29975 ;
  assign n29977 = n29976 ^ n29972 ;
  assign n30064 = n29977 ^ n28013 ;
  assign n30065 = n30064 ^ x502 ;
  assign n30248 = n30139 ^ n30065 ;
  assign n30249 = ~n30247 & ~n30248 ;
  assign n30140 = n30139 ^ n30064 ;
  assign n30141 = n30065 & ~n30140 ;
  assign n30142 = n30141 ^ x502 ;
  assign n29895 = n29811 ^ n29246 ;
  assign n29896 = n29895 ^ n28398 ;
  assign n29978 = ~n29896 & n29977 ;
  assign n29611 = n29610 ^ n29246 ;
  assign n29799 = n29611 & n29798 ;
  assign n29800 = n29799 ^ n29246 ;
  assign n29608 = n29456 ^ n29455 ;
  assign n29609 = n29608 ^ n29145 ;
  assign n29891 = n29800 ^ n29609 ;
  assign n29892 = n29891 ^ n29145 ;
  assign n29893 = n29892 ^ n29142 ;
  assign n29894 = n29893 ^ n28013 ;
  assign n29979 = n29978 ^ n29894 ;
  assign n30062 = n29979 ^ n28023 ;
  assign n30063 = n30062 ^ x501 ;
  assign n30250 = n30142 ^ n30063 ;
  assign n30251 = ~n30249 & n30250 ;
  assign n30143 = n30142 ^ n30062 ;
  assign n30144 = n30063 & ~n30143 ;
  assign n30145 = n30144 ^ x501 ;
  assign n29980 = n29892 ^ n28424 ;
  assign n29981 = ~n29979 & ~n29980 ;
  assign n29804 = n29458 ^ n29457 ;
  assign n29805 = n29804 ^ n29269 ;
  assign n29801 = n29800 ^ n29608 ;
  assign n29802 = n29609 & n29801 ;
  assign n29803 = n29802 ^ n29145 ;
  assign n29806 = n29805 ^ n29803 ;
  assign n29888 = n29806 ^ n29269 ;
  assign n29889 = n29888 ^ n29262 ;
  assign n29890 = n29889 ^ n28023 ;
  assign n29982 = n29981 ^ n29890 ;
  assign n30060 = n29982 ^ n27909 ;
  assign n30061 = n30060 ^ x500 ;
  assign n30252 = n30145 ^ n30061 ;
  assign n30253 = n30251 & ~n30252 ;
  assign n30146 = n30145 ^ n30060 ;
  assign n30147 = ~n30061 & n30146 ;
  assign n30148 = n30147 ^ x500 ;
  assign n29828 = n29460 ^ n29459 ;
  assign n29883 = n29828 ^ n29282 ;
  assign n29825 = n29804 ^ n29803 ;
  assign n29826 = n29805 & ~n29825 ;
  assign n29827 = n29826 ^ n29269 ;
  assign n29884 = n29883 ^ n29827 ;
  assign n29885 = n29884 ^ n29282 ;
  assign n29886 = n29885 ^ n29275 ;
  assign n29984 = n29886 ^ n27909 ;
  assign n29983 = n29889 ^ n29886 ;
  assign n29985 = n29984 ^ n29983 ;
  assign n29986 = n29982 & ~n29985 ;
  assign n29987 = n29986 ^ n29984 ;
  assign n30058 = n29987 ^ n27906 ;
  assign n30059 = n30058 ^ x499 ;
  assign n30254 = n30148 ^ n30059 ;
  assign n30255 = n30253 & n30254 ;
  assign n30149 = n30148 ^ n30058 ;
  assign n30150 = n30059 & ~n30149 ;
  assign n30151 = n30150 ^ x499 ;
  assign n29887 = n29886 ^ n27906 ;
  assign n29988 = n29887 & n29987 ;
  assign n29989 = n29988 ^ n27906 ;
  assign n30055 = n29989 ^ n27903 ;
  assign n29829 = n29828 ^ n29827 ;
  assign n29830 = n29462 ^ n29461 ;
  assign n29831 = n29830 ^ n29282 ;
  assign n29832 = n29831 ^ n29827 ;
  assign n29833 = n29832 ^ n29830 ;
  assign n29834 = n29829 & n29833 ;
  assign n29835 = n29834 ^ n29831 ;
  assign n29990 = n29835 ^ n29286 ;
  assign n30056 = n30055 ^ n29990 ;
  assign n30057 = n30056 ^ x498 ;
  assign n30256 = n30151 ^ n30057 ;
  assign n30257 = ~n30255 & ~n30256 ;
  assign n30152 = n30151 ^ n30056 ;
  assign n30153 = n30057 & ~n30152 ;
  assign n30154 = n30153 ^ x498 ;
  assign n29991 = n29990 ^ n29989 ;
  assign n29823 = n29464 ^ n29463 ;
  assign n29837 = n29823 ^ n29293 ;
  assign n29836 = n29830 ^ n29823 ;
  assign n29838 = n29837 ^ n29836 ;
  assign n29839 = ~n29835 & ~n29838 ;
  assign n29840 = n29839 ^ n29837 ;
  assign n29881 = n29840 ^ n29424 ;
  assign n29992 = n29881 ^ n27903 ;
  assign n29993 = n29992 ^ n29989 ;
  assign n29994 = n29993 ^ n29881 ;
  assign n29995 = n29991 & n29994 ;
  assign n29996 = n29995 ^ n29992 ;
  assign n30053 = n29996 ^ n27900 ;
  assign n30054 = n30053 ^ x497 ;
  assign n30258 = n30154 ^ n30054 ;
  assign n30259 = ~n30257 & ~n30258 ;
  assign n29822 = n29466 ^ n29465 ;
  assign n29999 = n29822 ^ n29495 ;
  assign n29824 = n29823 ^ n29430 ;
  assign n29841 = ~n29824 & ~n29840 ;
  assign n29842 = n29841 ^ n29430 ;
  assign n30000 = n29999 ^ n29842 ;
  assign n30001 = n30000 ^ n29495 ;
  assign n30002 = n30001 ^ n28766 ;
  assign n30159 = n30002 ^ n28047 ;
  assign n29882 = n29881 ^ n27900 ;
  assign n29997 = n29882 & n29996 ;
  assign n29998 = n29997 ^ n27900 ;
  assign n30160 = n30159 ^ n29998 ;
  assign n30155 = n30154 ^ n30053 ;
  assign n30156 = ~n30054 & n30155 ;
  assign n30157 = n30156 ^ x497 ;
  assign n30158 = n30157 ^ x496 ;
  assign n30218 = n30160 ^ n30158 ;
  assign n30290 = n30259 ^ n30218 ;
  assign n30293 = n30292 ^ n30290 ;
  assign n30297 = n29732 ^ n29724 ;
  assign n30296 = n30258 ^ n30257 ;
  assign n30298 = n30297 ^ n30296 ;
  assign n30300 = n29729 ^ n29148 ;
  assign n30301 = n30300 ^ n29725 ;
  assign n30299 = n30256 ^ n30255 ;
  assign n30302 = n30301 ^ n30299 ;
  assign n30304 = n29561 ^ n29173 ;
  assign n30305 = n30304 ^ n29582 ;
  assign n30303 = n30254 ^ n30253 ;
  assign n30306 = n30305 ^ n30303 ;
  assign n30310 = n30252 ^ n30251 ;
  assign n30307 = n29516 ^ n29167 ;
  assign n30308 = n30307 ^ n29539 ;
  assign n30311 = n30310 ^ n30308 ;
  assign n30313 = n29504 ^ n29161 ;
  assign n30314 = n30313 ^ n29512 ;
  assign n30312 = n30250 ^ n30249 ;
  assign n30315 = n30314 ^ n30312 ;
  assign n30317 = n30246 ^ n30219 ;
  assign n30318 = n29545 ^ n29033 ;
  assign n30319 = ~n30317 & ~n30318 ;
  assign n30324 = n30319 ^ n30312 ;
  assign n30316 = n30248 ^ n30247 ;
  assign n30320 = n30319 ^ n30316 ;
  assign n30321 = n29509 ^ n29508 ;
  assign n30322 = n30321 ^ n30316 ;
  assign n30323 = ~n30320 & ~n30322 ;
  assign n30325 = n30324 ^ n30323 ;
  assign n30326 = ~n30315 & n30325 ;
  assign n30327 = n30326 ^ n30314 ;
  assign n30328 = n30327 ^ n30308 ;
  assign n30329 = ~n30311 & n30328 ;
  assign n30309 = n30308 ^ n30303 ;
  assign n30330 = n30329 ^ n30309 ;
  assign n30331 = ~n30306 & ~n30330 ;
  assign n30332 = n30331 ^ n30305 ;
  assign n30333 = n30332 ^ n30299 ;
  assign n30334 = n30302 & ~n30333 ;
  assign n30335 = n30334 ^ n30301 ;
  assign n30336 = n30335 ^ n30296 ;
  assign n30337 = n30298 & n30336 ;
  assign n30338 = n30337 ^ n30297 ;
  assign n30260 = n30218 & ~n30259 ;
  assign n30003 = n30002 ^ n29998 ;
  assign n29843 = n29842 ^ n29822 ;
  assign n29844 = n29842 ^ n29495 ;
  assign n29845 = ~n29843 & n29844 ;
  assign n29846 = n29845 ^ n29495 ;
  assign n29820 = n29467 ^ n29442 ;
  assign n29821 = n29820 ^ n29528 ;
  assign n30004 = n29846 ^ n29821 ;
  assign n30005 = n30004 ^ n29528 ;
  assign n30006 = n30005 ^ n28818 ;
  assign n30007 = n30006 ^ n28047 ;
  assign n30008 = n30007 ^ n29998 ;
  assign n30009 = n30008 ^ n30006 ;
  assign n30010 = ~n30003 & ~n30009 ;
  assign n30011 = n30010 ^ n30007 ;
  assign n30052 = n30011 ^ n28210 ;
  assign n30216 = n30052 ^ x511 ;
  assign n30161 = n30160 ^ n30157 ;
  assign n30162 = n30158 & n30161 ;
  assign n30163 = n30162 ^ x496 ;
  assign n30217 = n30216 ^ n30163 ;
  assign n30288 = n30260 ^ n30217 ;
  assign n30294 = n30292 ^ n30288 ;
  assign n30295 = n30294 ^ n30288 ;
  assign n30339 = n30338 ^ n30295 ;
  assign n30340 = n30293 & n30339 ;
  assign n30341 = n30340 ^ n30294 ;
  assign n30287 = n29738 ^ n29720 ;
  assign n30457 = n30341 ^ n30287 ;
  assign n30405 = n30317 ^ n29033 ;
  assign n30406 = n30405 ^ x71 ;
  assign n30478 = n30321 ^ n30319 ;
  assign n30479 = n30478 ^ n30316 ;
  assign n30480 = n30479 ^ n29510 ;
  assign n30476 = n29034 & n30405 ;
  assign n30477 = n30476 ^ n29036 ;
  assign n30685 = n30480 ^ n30477 ;
  assign n30683 = x71 & ~n30405 ;
  assign n30684 = n30683 ^ x70 ;
  assign n30859 = n30685 ^ n30684 ;
  assign n30860 = ~n30406 & n30859 ;
  assign n30481 = n30480 ^ n30476 ;
  assign n30482 = n30477 & ~n30481 ;
  assign n30483 = n30482 ^ n29036 ;
  assign n30681 = n30483 ^ n29031 ;
  assign n30474 = n30325 ^ n30314 ;
  assign n30475 = n30474 ^ n29513 ;
  assign n30682 = n30681 ^ n30475 ;
  assign n30861 = n30682 ^ x69 ;
  assign n30686 = n30685 ^ n30683 ;
  assign n30687 = n30684 & ~n30686 ;
  assign n30688 = n30687 ^ x70 ;
  assign n30862 = n30861 ^ n30688 ;
  assign n30863 = ~n30860 & n30862 ;
  assign n30689 = n30688 ^ n30682 ;
  assign n30484 = n30483 ^ n30475 ;
  assign n30471 = n30327 ^ n30311 ;
  assign n30472 = n30471 ^ n29540 ;
  assign n30485 = n30472 ^ n29031 ;
  assign n30486 = n30485 ^ n30472 ;
  assign n30487 = n30486 ^ n30475 ;
  assign n30488 = ~n30484 & ~n30487 ;
  assign n30489 = n30488 ^ n30485 ;
  assign n30690 = n30489 ^ n29026 ;
  assign n30691 = n30690 ^ x69 ;
  assign n30692 = n30691 ^ n30682 ;
  assign n30693 = n30692 ^ n30690 ;
  assign n30694 = n30689 & ~n30693 ;
  assign n30695 = n30694 ^ n30691 ;
  assign n30864 = n30695 ^ x68 ;
  assign n30865 = ~n30863 & n30864 ;
  assign n30473 = n30472 ^ n29026 ;
  assign n30490 = ~n30473 & n30489 ;
  assign n30491 = n30490 ^ n29026 ;
  assign n30696 = n30491 ^ n29049 ;
  assign n30468 = n30330 ^ n30305 ;
  assign n30469 = n30468 ^ n29583 ;
  assign n30697 = n30696 ^ n30469 ;
  assign n30699 = n30697 ^ x68 ;
  assign n30698 = n30697 ^ n30690 ;
  assign n30700 = n30699 ^ n30698 ;
  assign n30701 = ~n30695 & n30700 ;
  assign n30702 = n30701 ^ n30699 ;
  assign n30866 = n30702 ^ x67 ;
  assign n30867 = n30865 & ~n30866 ;
  assign n30470 = n30469 ^ n29049 ;
  assign n30492 = n30491 ^ n30469 ;
  assign n30493 = n30470 & n30492 ;
  assign n30494 = n30493 ^ n29049 ;
  assign n30465 = n30332 ^ n30302 ;
  assign n30466 = n30465 ^ n29730 ;
  assign n30467 = n30466 ^ n29052 ;
  assign n30679 = n30494 ^ n30467 ;
  assign n30704 = n30679 ^ x67 ;
  assign n30703 = n30697 ^ n30679 ;
  assign n30705 = n30704 ^ n30703 ;
  assign n30706 = n30702 & ~n30705 ;
  assign n30707 = n30706 ^ n30704 ;
  assign n30868 = n30707 ^ x66 ;
  assign n30869 = ~n30867 & ~n30868 ;
  assign n30495 = n30494 ^ n30466 ;
  assign n30496 = n30467 & n30495 ;
  assign n30497 = n30496 ^ n29052 ;
  assign n30710 = n30497 ^ n29060 ;
  assign n30462 = n30335 ^ n30298 ;
  assign n30463 = n30462 ^ n29733 ;
  assign n30711 = n30710 ^ n30463 ;
  assign n30870 = n30711 ^ x65 ;
  assign n30680 = n30679 ^ x66 ;
  assign n30708 = n30680 & ~n30707 ;
  assign n30709 = n30708 ^ x66 ;
  assign n30871 = n30870 ^ n30709 ;
  assign n30872 = n30869 & ~n30871 ;
  assign n30712 = n30711 ^ n30709 ;
  assign n30464 = n30463 ^ n29060 ;
  assign n30498 = n30497 ^ n30463 ;
  assign n30499 = ~n30464 & n30498 ;
  assign n30500 = n30499 ^ n29060 ;
  assign n30713 = n30500 ^ n29068 ;
  assign n30460 = n30338 ^ n30293 ;
  assign n30461 = n30460 ^ n29736 ;
  assign n30714 = n30713 ^ n30461 ;
  assign n30715 = n30714 ^ x65 ;
  assign n30716 = n30715 ^ n30709 ;
  assign n30717 = n30716 ^ n30714 ;
  assign n30718 = ~n30712 & n30717 ;
  assign n30719 = n30718 ^ n30715 ;
  assign n30873 = n30719 ^ x64 ;
  assign n30874 = ~n30872 & ~n30873 ;
  assign n30501 = n30500 ^ n30461 ;
  assign n30458 = n30457 ^ n29739 ;
  assign n30502 = n30458 ^ n29068 ;
  assign n30503 = n30502 ^ n30458 ;
  assign n30504 = n30503 ^ n30461 ;
  assign n30505 = ~n30501 & n30504 ;
  assign n30506 = n30505 ^ n30502 ;
  assign n30677 = n30506 ^ n29076 ;
  assign n30721 = n30677 ^ x64 ;
  assign n30720 = n30714 ^ n30677 ;
  assign n30722 = n30721 ^ n30720 ;
  assign n30723 = n30719 & ~n30722 ;
  assign n30724 = n30723 ^ n30721 ;
  assign n30875 = n30724 ^ x79 ;
  assign n30876 = n30874 & ~n30875 ;
  assign n30678 = n30677 ^ x79 ;
  assign n30725 = ~n30678 & n30724 ;
  assign n30726 = n30725 ^ x79 ;
  assign n30289 = n30288 ^ n30287 ;
  assign n30342 = n30289 & ~n30341 ;
  assign n30343 = n30342 ^ n30288 ;
  assign n30284 = n29718 ^ n29201 ;
  assign n30285 = n30284 ^ n29741 ;
  assign n30261 = n30217 & n30260 ;
  assign n30164 = n30163 ^ n30052 ;
  assign n30165 = n30163 ^ x511 ;
  assign n30166 = n30164 & n30165 ;
  assign n30167 = n30166 ^ x511 ;
  assign n30214 = n30167 ^ x510 ;
  assign n29819 = n29469 ^ n29468 ;
  assign n30012 = n29819 ^ n29576 ;
  assign n29847 = n29846 ^ n29820 ;
  assign n29848 = n29821 & n29847 ;
  assign n29849 = n29848 ^ n29528 ;
  assign n30013 = n30012 ^ n29849 ;
  assign n30016 = n30013 ^ n28210 ;
  assign n30017 = n30016 ^ n29574 ;
  assign n30014 = n30013 ^ n30006 ;
  assign n30015 = n30014 ^ n29574 ;
  assign n30018 = n30017 ^ n30015 ;
  assign n30019 = ~n30011 & n30018 ;
  assign n30020 = n30019 ^ n30017 ;
  assign n30050 = n30020 ^ n28225 ;
  assign n30215 = n30214 ^ n30050 ;
  assign n30283 = n30261 ^ n30215 ;
  assign n30286 = n30285 ^ n30283 ;
  assign n30510 = n30343 ^ n30286 ;
  assign n30511 = n30510 ^ n29742 ;
  assign n30459 = n30458 ^ n29076 ;
  assign n30507 = n30459 & ~n30506 ;
  assign n30508 = n30507 ^ n29076 ;
  assign n30509 = n30508 ^ n29084 ;
  assign n30675 = n30511 ^ n30509 ;
  assign n30676 = n30675 ^ x78 ;
  assign n30858 = n30726 ^ n30676 ;
  assign n30926 = n30876 ^ n30858 ;
  assign n30925 = n30405 ^ n29545 ;
  assign n31026 = n30926 ^ n30925 ;
  assign n31027 = ~n30318 & n31026 ;
  assign n31037 = n31027 ^ n30925 ;
  assign n31038 = n29505 & ~n31037 ;
  assign n30927 = n30925 & ~n30926 ;
  assign n30877 = ~n30858 & ~n30876 ;
  assign n30344 = n30343 ^ n30285 ;
  assign n30345 = ~n30286 & ~n30344 ;
  assign n30346 = n30345 ^ n30343 ;
  assign n30279 = n29767 ^ n29207 ;
  assign n30262 = ~n30215 & n30261 ;
  assign n30021 = n30013 ^ n29574 ;
  assign n30022 = n30021 ^ n28225 ;
  assign n30023 = ~n30020 & ~n30022 ;
  assign n30024 = n30023 ^ n28225 ;
  assign n29850 = n29849 ^ n29819 ;
  assign n29817 = n29471 ^ n29470 ;
  assign n29851 = n29817 ^ n29576 ;
  assign n29852 = n29851 ^ n29819 ;
  assign n29853 = n29852 ^ n29817 ;
  assign n29854 = ~n29850 & ~n29853 ;
  assign n29855 = n29854 ^ n29851 ;
  assign n29879 = n29855 ^ n29618 ;
  assign n29880 = n29879 ^ n28378 ;
  assign n30172 = n30024 ^ n29880 ;
  assign n30051 = n30050 ^ x510 ;
  assign n30168 = n30167 ^ n30050 ;
  assign n30169 = n30051 & ~n30168 ;
  assign n30170 = n30169 ^ x510 ;
  assign n30171 = n30170 ^ x509 ;
  assign n30213 = n30172 ^ n30171 ;
  assign n30278 = n30262 ^ n30213 ;
  assign n30280 = n30279 ^ n30278 ;
  assign n30455 = n30346 ^ n30280 ;
  assign n30456 = n30455 ^ n29767 ;
  assign n30731 = n30456 ^ n29092 ;
  assign n30512 = n30511 ^ n30508 ;
  assign n30513 = ~n30509 & ~n30512 ;
  assign n30514 = n30513 ^ n29084 ;
  assign n30732 = n30731 ^ n30514 ;
  assign n30727 = n30726 ^ n30675 ;
  assign n30728 = n30676 & ~n30727 ;
  assign n30729 = n30728 ^ x78 ;
  assign n30730 = n30729 ^ x77 ;
  assign n30857 = n30732 ^ n30730 ;
  assign n30924 = n30877 ^ n30857 ;
  assign n30928 = n30927 ^ n30924 ;
  assign n31034 = n30928 ^ n30479 ;
  assign n31035 = ~n30321 & n31034 ;
  assign n31036 = n31035 ^ n30479 ;
  assign n31039 = n31038 ^ n31036 ;
  assign n31040 = n31039 ^ n29154 ;
  assign n31025 = n30317 ^ n29506 ;
  assign n31028 = n31027 ^ n31025 ;
  assign n31032 = x7 & ~n31028 ;
  assign n31033 = n31032 ^ x6 ;
  assign n31586 = n31040 ^ n31033 ;
  assign n30263 = n30213 & n30262 ;
  assign n29816 = n29474 ^ n29472 ;
  assign n30029 = n29816 ^ n29649 ;
  assign n29818 = n29817 ^ n29638 ;
  assign n29856 = ~n29818 & ~n29855 ;
  assign n29857 = n29856 ^ n29638 ;
  assign n30030 = n30029 ^ n29857 ;
  assign n30031 = n30030 ^ n29649 ;
  assign n30032 = n30031 ^ n28839 ;
  assign n30025 = n30024 ^ n29879 ;
  assign n30026 = ~n29880 & ~n30025 ;
  assign n30027 = n30026 ^ n28378 ;
  assign n30028 = n30027 ^ n28409 ;
  assign n30177 = n30032 ^ n30028 ;
  assign n30173 = n30172 ^ n30170 ;
  assign n30174 = n30171 & n30173 ;
  assign n30175 = n30174 ^ x509 ;
  assign n30176 = n30175 ^ x508 ;
  assign n30212 = n30177 ^ n30176 ;
  assign n30276 = n30263 ^ n30212 ;
  assign n30281 = n30279 ^ n30276 ;
  assign n30282 = n30281 ^ n30276 ;
  assign n30347 = n30346 ^ n30282 ;
  assign n30348 = n30280 & n30347 ;
  assign n30349 = n30348 ^ n30281 ;
  assign n30275 = n29772 ^ n29213 ;
  assign n30452 = n30349 ^ n30275 ;
  assign n30453 = n30452 ^ n29772 ;
  assign n30454 = n30453 ^ n29100 ;
  assign n30515 = n30514 ^ n30456 ;
  assign n30516 = n30514 ^ n29092 ;
  assign n30517 = n30515 & n30516 ;
  assign n30518 = n30517 ^ n29092 ;
  assign n30519 = n30518 ^ n30453 ;
  assign n30520 = ~n30454 & ~n30519 ;
  assign n30521 = n30520 ^ n29100 ;
  assign n30264 = ~n30212 & n30263 ;
  assign n30033 = n30032 ^ n30027 ;
  assign n30034 = ~n30028 & ~n30033 ;
  assign n30035 = n30034 ^ n28409 ;
  assign n30048 = n30035 ^ n28643 ;
  assign n29862 = n29476 ^ n29475 ;
  assign n29875 = n29862 ^ n29635 ;
  assign n29858 = n29857 ^ n29816 ;
  assign n29859 = n29857 ^ n29649 ;
  assign n29860 = ~n29858 & n29859 ;
  assign n29861 = n29860 ^ n29649 ;
  assign n29876 = n29875 ^ n29861 ;
  assign n29877 = n29876 ^ n29635 ;
  assign n29878 = n29877 ^ n29632 ;
  assign n30049 = n30048 ^ n29878 ;
  assign n30210 = n30049 ^ x507 ;
  assign n30178 = n30177 ^ n30175 ;
  assign n30179 = n30176 & ~n30178 ;
  assign n30180 = n30179 ^ x508 ;
  assign n30211 = n30210 ^ n30180 ;
  assign n30274 = n30264 ^ n30211 ;
  assign n30449 = n30274 ^ n29950 ;
  assign n30277 = n30276 ^ n30275 ;
  assign n30350 = n30277 & ~n30349 ;
  assign n30351 = n30350 ^ n30276 ;
  assign n30450 = n30449 ^ n30351 ;
  assign n30451 = n30450 ^ n29951 ;
  assign n30522 = n30521 ^ n30451 ;
  assign n30523 = n30521 ^ n29107 ;
  assign n30524 = n30522 & n30523 ;
  assign n30525 = n30524 ^ n29107 ;
  assign n30744 = n30525 ^ n28624 ;
  assign n30352 = n30351 ^ n30274 ;
  assign n30265 = ~n30211 & n30264 ;
  assign n30181 = n30180 ^ n30049 ;
  assign n30182 = n30180 ^ x507 ;
  assign n30183 = ~n30181 & n30182 ;
  assign n30184 = n30183 ^ x507 ;
  assign n30036 = n30035 ^ n29878 ;
  assign n29863 = n29862 ^ n29861 ;
  assign n29814 = n29478 ^ n29477 ;
  assign n29864 = n29814 ^ n29635 ;
  assign n29865 = n29864 ^ n29814 ;
  assign n29866 = n29865 ^ n29861 ;
  assign n29867 = n29863 & n29866 ;
  assign n29868 = n29867 ^ n29864 ;
  assign n29873 = n29868 ^ n28854 ;
  assign n30037 = n29873 ^ n28643 ;
  assign n30038 = n30037 ^ n29878 ;
  assign n30039 = n30038 ^ n29873 ;
  assign n30040 = ~n30036 & n30039 ;
  assign n30041 = n30040 ^ n30037 ;
  assign n30046 = n30041 ^ n28662 ;
  assign n30047 = n30046 ^ x506 ;
  assign n30209 = n30184 ^ n30047 ;
  assign n30272 = n30265 ^ n30209 ;
  assign n30353 = n30272 ^ n29950 ;
  assign n30354 = n30353 ^ n30274 ;
  assign n30355 = n30354 ^ n30272 ;
  assign n30356 = ~n30352 & n30355 ;
  assign n30357 = n30356 ^ n30353 ;
  assign n30446 = n30357 ^ n29904 ;
  assign n30447 = n30446 ^ n29905 ;
  assign n30745 = n30744 ^ n30447 ;
  assign n30670 = n30451 ^ n29107 ;
  assign n30671 = n30670 ^ n30521 ;
  assign n30672 = n30671 ^ x75 ;
  assign n30733 = n30732 ^ n30729 ;
  assign n30734 = n30730 & n30733 ;
  assign n30735 = n30734 ^ x77 ;
  assign n30673 = n30518 ^ n29100 ;
  assign n30674 = n30673 ^ n30453 ;
  assign n30736 = n30735 ^ n30674 ;
  assign n30737 = n30735 ^ x76 ;
  assign n30738 = n30736 & n30737 ;
  assign n30739 = n30738 ^ x76 ;
  assign n30740 = n30739 ^ n30671 ;
  assign n30741 = n30672 & ~n30740 ;
  assign n30742 = n30741 ^ x75 ;
  assign n30743 = n30742 ^ x74 ;
  assign n30853 = n30745 ^ n30743 ;
  assign n30854 = n30739 ^ n30672 ;
  assign n30855 = n30674 ^ x76 ;
  assign n30856 = n30855 ^ n30735 ;
  assign n30878 = n30857 & n30877 ;
  assign n30879 = ~n30856 & ~n30878 ;
  assign n30880 = ~n30854 & ~n30879 ;
  assign n30881 = n30853 & ~n30880 ;
  assign n30273 = n30272 ^ n29904 ;
  assign n30358 = n30273 & n30357 ;
  assign n30359 = n30358 ^ n29904 ;
  assign n30443 = n30359 ^ n29900 ;
  assign n30266 = n30209 & ~n30265 ;
  assign n29874 = n29873 ^ n28662 ;
  assign n30042 = n29874 & n30041 ;
  assign n30043 = n30042 ^ n28662 ;
  assign n30044 = n30043 ^ n28681 ;
  assign n29815 = n29814 ^ n29685 ;
  assign n29869 = n29815 & ~n29868 ;
  assign n29870 = n29869 ^ n29685 ;
  assign n29813 = n29480 ^ n29479 ;
  assign n29871 = n29870 ^ n29813 ;
  assign n29872 = n29871 ^ n29703 ;
  assign n30045 = n30044 ^ n29872 ;
  assign n30207 = n30045 ^ x505 ;
  assign n30185 = n30184 ^ n30046 ;
  assign n30186 = n30047 & ~n30185 ;
  assign n30187 = n30186 ^ x506 ;
  assign n30208 = n30207 ^ n30187 ;
  assign n30271 = n30266 ^ n30208 ;
  assign n30444 = n30443 ^ n30271 ;
  assign n30445 = n30444 ^ n29901 ;
  assign n30668 = n30445 ^ n28621 ;
  assign n30448 = n30447 ^ n28624 ;
  assign n30526 = n30525 ^ n30447 ;
  assign n30527 = ~n30448 & ~n30526 ;
  assign n30528 = n30527 ^ n28624 ;
  assign n30669 = n30668 ^ n30528 ;
  assign n30851 = n30669 ^ x73 ;
  assign n30746 = n30745 ^ n30742 ;
  assign n30747 = n30743 & ~n30746 ;
  assign n30748 = n30747 ^ x74 ;
  assign n30852 = n30851 ^ n30748 ;
  assign n30945 = n30881 ^ n30852 ;
  assign n30921 = n30880 ^ n30853 ;
  assign n30922 = n30921 ^ n30468 ;
  assign n30929 = n30924 ^ n30479 ;
  assign n30930 = n30928 & ~n30929 ;
  assign n30931 = n30930 ^ n30479 ;
  assign n30932 = n30931 ^ n30474 ;
  assign n30933 = n30878 ^ n30856 ;
  assign n30934 = n30933 ^ n30931 ;
  assign n30935 = ~n30932 & ~n30934 ;
  assign n30936 = n30935 ^ n30474 ;
  assign n30923 = n30879 ^ n30854 ;
  assign n30937 = n30936 ^ n30923 ;
  assign n30938 = n30921 ^ n30471 ;
  assign n30939 = n30938 ^ n30923 ;
  assign n30940 = n30939 ^ n30921 ;
  assign n30941 = ~n30937 & n30940 ;
  assign n30942 = n30941 ^ n30938 ;
  assign n30943 = n30922 & ~n30942 ;
  assign n30944 = n30943 ^ n30468 ;
  assign n30946 = n30945 ^ n30944 ;
  assign n30882 = n30852 & ~n30881 ;
  assign n30749 = n30748 ^ n30669 ;
  assign n30750 = n30748 ^ x73 ;
  assign n30751 = n30749 & n30750 ;
  assign n30752 = n30751 ^ x73 ;
  assign n30529 = n30528 ^ n30445 ;
  assign n30530 = n30528 ^ n28621 ;
  assign n30531 = ~n30529 & ~n30530 ;
  assign n30532 = n30531 ^ n28621 ;
  assign n30665 = n30532 ^ n29128 ;
  assign n30360 = n30359 ^ n30271 ;
  assign n30269 = n29790 ^ n29236 ;
  assign n30361 = n30269 ^ n29900 ;
  assign n30362 = n30361 ^ n30271 ;
  assign n30363 = n30362 ^ n30269 ;
  assign n30364 = n30360 & ~n30363 ;
  assign n30365 = n30364 ^ n30361 ;
  assign n30267 = n30208 & n30266 ;
  assign n30203 = n30043 ^ n29872 ;
  assign n30204 = ~n30044 & ~n30203 ;
  assign n30194 = n29813 ^ n29709 ;
  assign n30195 = n29871 & ~n30194 ;
  assign n30191 = n29482 ^ n29481 ;
  assign n30192 = n30191 ^ n29751 ;
  assign n30193 = n30192 ^ n29813 ;
  assign n30196 = n30195 ^ n30193 ;
  assign n30197 = n30196 ^ n29751 ;
  assign n30198 = n30197 ^ n28877 ;
  assign n30199 = n30198 ^ n28681 ;
  assign n30200 = n30199 ^ n28722 ;
  assign n30201 = n30200 ^ x504 ;
  assign n30202 = n30201 ^ x505 ;
  assign n30205 = n30204 ^ n30202 ;
  assign n30188 = n30187 ^ n30045 ;
  assign n30189 = n30187 ^ x505 ;
  assign n30190 = ~n30188 & n30189 ;
  assign n30206 = n30205 ^ n30190 ;
  assign n30268 = n30267 ^ n30206 ;
  assign n30533 = n30365 ^ n30268 ;
  assign n30534 = n30533 ^ n29790 ;
  assign n30666 = n30665 ^ n30534 ;
  assign n30667 = n30666 ^ x72 ;
  assign n30850 = n30752 ^ n30667 ;
  assign n30947 = n30882 ^ n30850 ;
  assign n30948 = n30947 ^ n30465 ;
  assign n30949 = n30948 ^ n30944 ;
  assign n30950 = n30949 ^ n30947 ;
  assign n30951 = n30946 & n30950 ;
  assign n30952 = n30951 ^ n30948 ;
  assign n31030 = n30952 ^ n30462 ;
  assign n31029 = n31028 ^ x7 ;
  assign n31031 = n31030 ^ n31029 ;
  assign n31049 = n30933 ^ n30932 ;
  assign n31050 = n30314 & n31049 ;
  assign n31051 = n31050 ^ n30474 ;
  assign n31045 = n31036 ^ n29154 ;
  assign n31046 = n31039 & n31045 ;
  assign n31047 = n31046 ^ n29154 ;
  assign n31048 = n31047 ^ n29161 ;
  assign n31052 = n31051 ^ n31048 ;
  assign n31041 = n31040 ^ n31032 ;
  assign n31042 = n31033 & ~n31041 ;
  assign n31043 = n31042 ^ x6 ;
  assign n31044 = n31043 ^ x5 ;
  assign n31053 = n31052 ^ n31044 ;
  assign n31063 = n31051 ^ n31047 ;
  assign n31064 = n31051 ^ n29161 ;
  assign n31065 = n31063 & ~n31064 ;
  assign n31066 = n31065 ^ n29161 ;
  assign n31067 = n31066 ^ n29167 ;
  assign n31059 = n30936 ^ n30471 ;
  assign n31060 = n31059 ^ n30923 ;
  assign n31061 = n30308 & n31060 ;
  assign n31062 = n31061 ^ n30471 ;
  assign n31068 = n31067 ^ n31062 ;
  assign n31054 = n31052 ^ n31043 ;
  assign n31055 = n31052 ^ x5 ;
  assign n31056 = ~n31054 & n31055 ;
  assign n31057 = n31056 ^ x5 ;
  assign n31058 = n31057 ^ x4 ;
  assign n31069 = n31068 ^ n31058 ;
  assign n31070 = n31053 & n31069 ;
  assign n31080 = n31068 ^ n31057 ;
  assign n31081 = n31068 ^ x4 ;
  assign n31082 = ~n31080 & n31081 ;
  assign n31083 = n31082 ^ x4 ;
  assign n31084 = n31083 ^ x3 ;
  assign n31074 = n31062 ^ n29167 ;
  assign n31075 = n31066 ^ n31062 ;
  assign n31076 = ~n31074 & n31075 ;
  assign n31077 = n31076 ^ n29167 ;
  assign n31078 = n31077 ^ n29173 ;
  assign n31071 = n30942 ^ n30468 ;
  assign n31072 = ~n30305 & n31071 ;
  assign n31073 = n31072 ^ n30468 ;
  assign n31079 = n31078 ^ n31073 ;
  assign n31085 = n31084 ^ n31079 ;
  assign n31086 = n31070 & ~n31085 ;
  assign n31096 = n31079 ^ x3 ;
  assign n31097 = n31083 ^ n31079 ;
  assign n31098 = ~n31096 & n31097 ;
  assign n31099 = n31098 ^ x3 ;
  assign n31100 = n31099 ^ x2 ;
  assign n31092 = n31077 ^ n31073 ;
  assign n31093 = ~n31078 & n31092 ;
  assign n31094 = n31093 ^ n29173 ;
  assign n31087 = n30945 ^ n30465 ;
  assign n31088 = n31087 ^ n30944 ;
  assign n31089 = ~n30301 & ~n31088 ;
  assign n31090 = n31089 ^ n30465 ;
  assign n31091 = n31090 ^ n29148 ;
  assign n31095 = n31094 ^ n31091 ;
  assign n31101 = n31100 ^ n31095 ;
  assign n31102 = n31086 & ~n31101 ;
  assign n31112 = n31099 ^ n31095 ;
  assign n31113 = n31100 & n31112 ;
  assign n31114 = n31113 ^ x2 ;
  assign n31105 = n31094 ^ n31090 ;
  assign n31106 = n31094 ^ n29148 ;
  assign n31107 = ~n31105 & ~n31106 ;
  assign n31108 = n31107 ^ n29148 ;
  assign n31109 = n31108 ^ n29183 ;
  assign n31103 = n30297 & n31030 ;
  assign n31104 = n31103 ^ n30462 ;
  assign n31110 = n31109 ^ n31104 ;
  assign n31111 = n31110 ^ x1 ;
  assign n31115 = n31114 ^ n31111 ;
  assign n31116 = ~n31102 & ~n31115 ;
  assign n31127 = n31114 ^ n31110 ;
  assign n31128 = n31114 ^ x1 ;
  assign n31129 = ~n31127 & n31128 ;
  assign n31130 = n31129 ^ x1 ;
  assign n31131 = n31130 ^ x0 ;
  assign n31117 = n31108 ^ n31104 ;
  assign n30883 = n30850 & ~n30882 ;
  assign n30368 = n29589 ^ x487 ;
  assign n30539 = n30368 ^ n29967 ;
  assign n30270 = n30269 ^ n30268 ;
  assign n30366 = n30270 & ~n30365 ;
  assign n30367 = n30366 ^ n30269 ;
  assign n30540 = n30539 ^ n30367 ;
  assign n30541 = n30540 ^ n29968 ;
  assign n30663 = n30541 ^ n29125 ;
  assign n30535 = n30534 ^ n30532 ;
  assign n30536 = n30534 ^ n29128 ;
  assign n30537 = n30535 & ~n30536 ;
  assign n30538 = n30537 ^ n29128 ;
  assign n30664 = n30663 ^ n30538 ;
  assign n30848 = n30664 ^ x87 ;
  assign n30753 = n30752 ^ n30666 ;
  assign n30754 = n30667 & ~n30753 ;
  assign n30755 = n30754 ^ x72 ;
  assign n30849 = n30848 ^ n30755 ;
  assign n30919 = n30883 ^ n30849 ;
  assign n30954 = n30919 ^ n30462 ;
  assign n30953 = n30947 ^ n30919 ;
  assign n30955 = n30954 ^ n30953 ;
  assign n30956 = ~n30952 & n30955 ;
  assign n30957 = n30956 ^ n30954 ;
  assign n31118 = n30957 ^ n30460 ;
  assign n31119 = n30292 & n31118 ;
  assign n31120 = n31119 ^ n30460 ;
  assign n31121 = n31120 ^ n29183 ;
  assign n31122 = n31121 ^ n31120 ;
  assign n31123 = n31122 ^ n31108 ;
  assign n31124 = n31117 & n31123 ;
  assign n31125 = n31124 ^ n31121 ;
  assign n31126 = n31125 ^ n29189 ;
  assign n31132 = n31131 ^ n31126 ;
  assign n31133 = ~n31116 & ~n31132 ;
  assign n31134 = n31130 ^ n31126 ;
  assign n31147 = n31131 & n31134 ;
  assign n31139 = n31120 ^ n29189 ;
  assign n31140 = ~n31125 & n31139 ;
  assign n31141 = n31140 ^ n29189 ;
  assign n31142 = n31141 ^ n29195 ;
  assign n30884 = n30849 & n30883 ;
  assign n30542 = n30541 ^ n30538 ;
  assign n30369 = n30368 ^ n30367 ;
  assign n30372 = n30367 ^ n29967 ;
  assign n30373 = ~n30369 & n30372 ;
  assign n30370 = n29967 ^ n29811 ;
  assign n30374 = n30373 ^ n30370 ;
  assign n29810 = n29592 ^ n29591 ;
  assign n30440 = n30374 ^ n29810 ;
  assign n30441 = n30440 ^ n29895 ;
  assign n30543 = n30441 ^ n29125 ;
  assign n30544 = n30543 ^ n30441 ;
  assign n30545 = n30544 ^ n30538 ;
  assign n30546 = ~n30542 & ~n30545 ;
  assign n30547 = n30546 ^ n30543 ;
  assign n30760 = n30547 ^ n29139 ;
  assign n30846 = n30760 ^ x86 ;
  assign n30756 = n30755 ^ n30664 ;
  assign n30757 = n30755 ^ x87 ;
  assign n30758 = ~n30756 & n30757 ;
  assign n30759 = n30758 ^ x87 ;
  assign n30847 = n30846 ^ n30759 ;
  assign n30918 = n30884 ^ n30847 ;
  assign n31135 = n30918 ^ n30457 ;
  assign n30920 = n30919 ^ n30460 ;
  assign n30958 = n30920 & n30957 ;
  assign n30959 = n30958 ^ n30460 ;
  assign n31136 = n31135 ^ n30959 ;
  assign n31137 = ~n30287 & ~n31136 ;
  assign n31138 = n31137 ^ n30457 ;
  assign n31143 = n31142 ^ n31138 ;
  assign n31144 = n31143 ^ x0 ;
  assign n31148 = n31147 ^ n31144 ;
  assign n31149 = n31148 ^ x15 ;
  assign n31150 = n31133 & n31149 ;
  assign n31159 = n31143 ^ x15 ;
  assign n31160 = ~n31148 & n31159 ;
  assign n31161 = n31160 ^ x15 ;
  assign n31162 = n31161 ^ x14 ;
  assign n31154 = n31141 ^ n31138 ;
  assign n31155 = ~n31142 & ~n31154 ;
  assign n31156 = n31155 ^ n29195 ;
  assign n31157 = n31156 ^ n29201 ;
  assign n30960 = n30959 ^ n30918 ;
  assign n30961 = n30959 ^ n30457 ;
  assign n30962 = ~n30960 & n30961 ;
  assign n30963 = n30962 ^ n30457 ;
  assign n30885 = n30847 & n30884 ;
  assign n30761 = n30760 ^ n30759 ;
  assign n29808 = n29595 ^ x485 ;
  assign n29809 = n29808 ^ n29588 ;
  assign n30551 = n29891 ^ n29809 ;
  assign n29812 = n29811 ^ n29810 ;
  assign n30375 = n29812 & ~n30374 ;
  assign n30376 = n30375 ^ n29811 ;
  assign n30552 = n30551 ^ n30376 ;
  assign n30553 = n30552 ^ n29892 ;
  assign n30442 = n30441 ^ n29139 ;
  assign n30548 = n30442 & ~n30547 ;
  assign n30549 = n30548 ^ n29139 ;
  assign n30550 = n30549 ^ n29142 ;
  assign n30661 = n30553 ^ n30550 ;
  assign n30762 = n30661 ^ x86 ;
  assign n30763 = n30762 ^ n30661 ;
  assign n30764 = n30763 ^ n30759 ;
  assign n30765 = ~n30761 & n30764 ;
  assign n30766 = n30765 ^ n30762 ;
  assign n30845 = n30766 ^ x85 ;
  assign n30916 = n30885 ^ n30845 ;
  assign n30917 = n30916 ^ n30510 ;
  assign n31151 = n30963 ^ n30917 ;
  assign n31152 = n30285 & ~n31151 ;
  assign n31153 = n31152 ^ n30510 ;
  assign n31158 = n31157 ^ n31153 ;
  assign n31163 = n31162 ^ n31158 ;
  assign n31164 = ~n31150 & ~n31163 ;
  assign n31174 = n31161 ^ n31158 ;
  assign n31175 = n31162 & ~n31174 ;
  assign n31176 = n31175 ^ x14 ;
  assign n31168 = n31156 ^ n31153 ;
  assign n31169 = n31157 & ~n31168 ;
  assign n31170 = n31169 ^ n29201 ;
  assign n31171 = n31170 ^ n29207 ;
  assign n30886 = ~n30845 & ~n30885 ;
  assign n30377 = n30376 ^ n29809 ;
  assign n30378 = n30376 ^ n29891 ;
  assign n30379 = ~n30377 & n30378 ;
  assign n30380 = n30379 ^ n29891 ;
  assign n29807 = n29806 ^ n29606 ;
  assign n30438 = n30380 ^ n29807 ;
  assign n30439 = n30438 ^ n29888 ;
  assign n30769 = n30439 ^ n29262 ;
  assign n30554 = n30553 ^ n30549 ;
  assign n30555 = n30550 & ~n30554 ;
  assign n30556 = n30555 ^ n29142 ;
  assign n30770 = n30769 ^ n30556 ;
  assign n30843 = n30770 ^ x84 ;
  assign n30662 = n30661 ^ x85 ;
  assign n30767 = n30662 & ~n30766 ;
  assign n30768 = n30767 ^ x85 ;
  assign n30844 = n30843 ^ n30768 ;
  assign n30968 = n30886 ^ n30844 ;
  assign n30964 = n30963 ^ n30916 ;
  assign n30965 = n30917 & n30964 ;
  assign n30966 = n30965 ^ n30510 ;
  assign n30967 = n30966 ^ n30455 ;
  assign n31165 = n30968 ^ n30967 ;
  assign n31166 = ~n30279 & ~n31165 ;
  assign n31167 = n31166 ^ n30455 ;
  assign n31172 = n31171 ^ n31167 ;
  assign n31173 = n31172 ^ x13 ;
  assign n31177 = n31176 ^ n31173 ;
  assign n31178 = ~n31164 & ~n31177 ;
  assign n31183 = n31170 ^ n31167 ;
  assign n30887 = ~n30844 & n30886 ;
  assign n30771 = n30770 ^ n30768 ;
  assign n30557 = n30556 ^ n30439 ;
  assign n30558 = n30556 ^ n29262 ;
  assign n30559 = n30557 & ~n30558 ;
  assign n30560 = n30559 ^ n29262 ;
  assign n29607 = n29606 ^ n29605 ;
  assign n30434 = n29884 ^ n29607 ;
  assign n30381 = n30380 ^ n29806 ;
  assign n30382 = n29807 & n30381 ;
  assign n30383 = n30382 ^ n29606 ;
  assign n30435 = n30434 ^ n30383 ;
  assign n30436 = n30435 ^ n29885 ;
  assign n30437 = n30436 ^ n29275 ;
  assign n30772 = n30560 ^ n30437 ;
  assign n30773 = n30772 ^ x84 ;
  assign n30774 = n30773 ^ n30768 ;
  assign n30775 = n30774 ^ n30772 ;
  assign n30776 = ~n30771 & n30775 ;
  assign n30777 = n30776 ^ n30773 ;
  assign n30842 = n30777 ^ x83 ;
  assign n30915 = n30887 ^ n30842 ;
  assign n31184 = n30915 ^ n30452 ;
  assign n30969 = n30968 ^ n30966 ;
  assign n30970 = n30967 & n30969 ;
  assign n30971 = n30970 ^ n30455 ;
  assign n31185 = n31184 ^ n30971 ;
  assign n31186 = n30275 & n31185 ;
  assign n31187 = n31186 ^ n30452 ;
  assign n31188 = n31187 ^ n29207 ;
  assign n31189 = n31188 ^ n31167 ;
  assign n31190 = n31189 ^ n31187 ;
  assign n31191 = ~n31183 & ~n31190 ;
  assign n31192 = n31191 ^ n31188 ;
  assign n31193 = n31192 ^ n29213 ;
  assign n31194 = n31193 ^ x12 ;
  assign n31179 = n31176 ^ n31172 ;
  assign n31180 = n31176 ^ x13 ;
  assign n31181 = n31179 & n31180 ;
  assign n31182 = n31181 ^ x13 ;
  assign n31195 = n31194 ^ n31182 ;
  assign n31196 = n31178 & n31195 ;
  assign n31204 = n31187 ^ n29213 ;
  assign n31205 = n31192 & ~n31204 ;
  assign n31206 = n31205 ^ n29213 ;
  assign n30972 = n30971 ^ n30915 ;
  assign n30973 = n30971 ^ n30452 ;
  assign n30974 = ~n30972 & n30973 ;
  assign n30975 = n30974 ^ n30452 ;
  assign n30888 = n30842 & ~n30887 ;
  assign n30391 = n30223 ^ n30221 ;
  assign n30388 = n29835 ^ n29293 ;
  assign n30431 = n30391 ^ n30388 ;
  assign n30384 = n30383 ^ n29607 ;
  assign n30385 = n30383 ^ n29884 ;
  assign n30386 = n30384 & ~n30385 ;
  assign n30387 = n30386 ^ n29884 ;
  assign n30432 = n30431 ^ n30387 ;
  assign n30433 = n30432 ^ n29835 ;
  assign n30778 = n30433 ^ n29286 ;
  assign n30561 = n30560 ^ n30436 ;
  assign n30562 = ~n30437 & ~n30561 ;
  assign n30563 = n30562 ^ n29275 ;
  assign n30779 = n30778 ^ n30563 ;
  assign n30781 = n30779 ^ x83 ;
  assign n30780 = n30779 ^ n30772 ;
  assign n30782 = n30781 ^ n30780 ;
  assign n30783 = ~n30777 & n30782 ;
  assign n30784 = n30783 ^ n30781 ;
  assign n30841 = n30784 ^ x82 ;
  assign n30913 = n30888 ^ n30841 ;
  assign n30914 = n30913 ^ n30450 ;
  assign n31200 = n30975 ^ n30914 ;
  assign n31201 = n29950 & ~n31200 ;
  assign n31202 = n31201 ^ n30450 ;
  assign n31203 = n31202 ^ n29219 ;
  assign n31207 = n31206 ^ n31203 ;
  assign n31208 = n31207 ^ x11 ;
  assign n31197 = n31193 ^ n31182 ;
  assign n31198 = n31194 & ~n31197 ;
  assign n31199 = n31198 ^ x12 ;
  assign n31209 = n31208 ^ n31199 ;
  assign n31210 = n31196 & n31209 ;
  assign n31211 = n31207 ^ n31199 ;
  assign n30889 = ~n30841 & ~n30888 ;
  assign n30564 = n30563 ^ n30433 ;
  assign n30565 = n30563 ^ n29286 ;
  assign n30566 = ~n30564 & n30565 ;
  assign n30567 = n30566 ^ n29286 ;
  assign n30658 = n30567 ^ n29424 ;
  assign n30398 = n30224 ^ n30220 ;
  assign n30389 = n30388 ^ n30387 ;
  assign n30394 = n30391 ^ n30387 ;
  assign n30395 = ~n30389 & ~n30394 ;
  assign n30390 = n29840 ^ n29430 ;
  assign n30392 = n30391 ^ n30390 ;
  assign n30396 = n30395 ^ n30392 ;
  assign n30428 = n30398 ^ n30396 ;
  assign n30429 = n30428 ^ n29840 ;
  assign n30659 = n30658 ^ n30429 ;
  assign n30786 = n30659 ^ x82 ;
  assign n30785 = n30779 ^ n30659 ;
  assign n30787 = n30786 ^ n30785 ;
  assign n30788 = ~n30784 & n30787 ;
  assign n30789 = n30788 ^ n30786 ;
  assign n30840 = n30789 ^ x81 ;
  assign n30979 = n30889 ^ n30840 ;
  assign n31216 = n30979 ^ n30446 ;
  assign n30976 = n30975 ^ n30913 ;
  assign n30977 = ~n30914 & ~n30976 ;
  assign n30978 = n30977 ^ n30450 ;
  assign n31217 = n31216 ^ n30978 ;
  assign n31218 = ~n29904 & ~n31217 ;
  assign n31219 = n31218 ^ n30446 ;
  assign n31220 = n31219 ^ n29225 ;
  assign n31212 = n31206 ^ n31202 ;
  assign n31213 = n31206 ^ n29219 ;
  assign n31214 = ~n31212 & ~n31213 ;
  assign n31215 = n31214 ^ n29219 ;
  assign n31221 = n31220 ^ n31215 ;
  assign n31222 = n31221 ^ x11 ;
  assign n31223 = n31222 ^ n31199 ;
  assign n31224 = n31223 ^ n31221 ;
  assign n31225 = ~n31211 & n31224 ;
  assign n31226 = n31225 ^ n31222 ;
  assign n31227 = n31226 ^ x10 ;
  assign n31228 = ~n31210 & n31227 ;
  assign n30980 = n30979 ^ n30978 ;
  assign n30890 = ~n30840 & ~n30889 ;
  assign n30430 = n30429 ^ n29424 ;
  assign n30568 = n30567 ^ n30429 ;
  assign n30569 = ~n30430 & n30568 ;
  assign n30570 = n30569 ^ n29424 ;
  assign n30656 = n30570 ^ n28766 ;
  assign n30397 = n30227 ^ n30225 ;
  assign n30400 = n30397 ^ n30390 ;
  assign n30399 = n30398 ^ n30397 ;
  assign n30401 = n30400 ^ n30399 ;
  assign n30402 = n30396 & ~n30401 ;
  assign n30403 = n30402 ^ n30400 ;
  assign n30404 = n30403 ^ n30000 ;
  assign n30427 = n30404 ^ n30001 ;
  assign n30657 = n30656 ^ n30427 ;
  assign n30838 = n30657 ^ x80 ;
  assign n30660 = n30659 ^ x81 ;
  assign n30790 = ~n30660 & n30789 ;
  assign n30791 = n30790 ^ x81 ;
  assign n30839 = n30838 ^ n30791 ;
  assign n30911 = n30890 ^ n30839 ;
  assign n30981 = n30911 ^ n30446 ;
  assign n30982 = n30981 ^ n30978 ;
  assign n30983 = n30982 ^ n30911 ;
  assign n30984 = ~n30980 & n30983 ;
  assign n30985 = n30984 ^ n30981 ;
  assign n31232 = n30985 ^ n30444 ;
  assign n31233 = ~n29900 & n31232 ;
  assign n31234 = n31233 ^ n30444 ;
  assign n31235 = n31234 ^ n29231 ;
  assign n31229 = n31219 ^ n31215 ;
  assign n31230 = ~n31220 & n31229 ;
  assign n31231 = n31230 ^ n29225 ;
  assign n31236 = n31235 ^ n31231 ;
  assign n31238 = n31236 ^ x10 ;
  assign n31237 = n31236 ^ n31221 ;
  assign n31239 = n31238 ^ n31237 ;
  assign n31240 = n31226 & ~n31239 ;
  assign n31241 = n31240 ^ n31238 ;
  assign n31242 = n31241 ^ x9 ;
  assign n31243 = ~n31228 & n31242 ;
  assign n31244 = n31234 ^ n31231 ;
  assign n30891 = ~n30839 & ~n30890 ;
  assign n30792 = n30791 ^ n30657 ;
  assign n30793 = n30791 ^ x80 ;
  assign n30794 = ~n30792 & n30793 ;
  assign n30795 = n30794 ^ x80 ;
  assign n30571 = n30570 ^ n30427 ;
  assign n30413 = n30229 ^ n30228 ;
  assign n30572 = n30413 ^ n30004 ;
  assign n30414 = n30397 ^ n30000 ;
  assign n30415 = ~n30403 & n30414 ;
  assign n30416 = n30415 ^ n30000 ;
  assign n30573 = n30572 ^ n30416 ;
  assign n30574 = n30573 ^ n30005 ;
  assign n30575 = n30574 ^ n28766 ;
  assign n30576 = n30575 ^ n30427 ;
  assign n30577 = n30576 ^ n30574 ;
  assign n30578 = ~n30571 & n30577 ;
  assign n30579 = n30578 ^ n30575 ;
  assign n30654 = n30579 ^ n28818 ;
  assign n30655 = n30654 ^ x95 ;
  assign n30837 = n30795 ^ n30655 ;
  assign n30910 = n30891 ^ n30837 ;
  assign n31245 = n30910 ^ n30533 ;
  assign n30912 = n30911 ^ n30444 ;
  assign n30986 = ~n30912 & n30985 ;
  assign n30987 = n30986 ^ n30444 ;
  assign n31246 = n31245 ^ n30987 ;
  assign n31247 = n30269 & n31246 ;
  assign n31248 = n31247 ^ n30533 ;
  assign n31249 = n31248 ^ n29231 ;
  assign n31250 = n31249 ^ n31231 ;
  assign n31251 = n31250 ^ n31248 ;
  assign n31252 = n31244 & ~n31251 ;
  assign n31253 = n31252 ^ n31249 ;
  assign n31254 = n31253 ^ n29236 ;
  assign n31256 = n31254 ^ x9 ;
  assign n31255 = n31254 ^ n31236 ;
  assign n31257 = n31256 ^ n31255 ;
  assign n31258 = ~n31241 & n31257 ;
  assign n31259 = n31258 ^ n31256 ;
  assign n31260 = n31259 ^ x8 ;
  assign n31261 = n31243 & n31260 ;
  assign n31266 = n31248 ^ n29236 ;
  assign n31267 = n31253 & ~n31266 ;
  assign n31268 = n31267 ^ n29236 ;
  assign n30988 = n30987 ^ n30910 ;
  assign n30989 = n30987 ^ n30533 ;
  assign n30990 = ~n30988 & ~n30989 ;
  assign n30991 = n30990 ^ n30533 ;
  assign n30892 = ~n30837 & ~n30891 ;
  assign n30581 = n30013 ^ n29576 ;
  assign n30417 = n30416 ^ n30413 ;
  assign n30418 = n30416 ^ n30004 ;
  assign n30419 = ~n30417 & n30418 ;
  assign n30420 = n30419 ^ n30004 ;
  assign n30411 = n30231 ^ n30230 ;
  assign n30412 = n30411 ^ n30013 ;
  assign n30580 = n30420 ^ n30412 ;
  assign n30582 = n30581 ^ n30580 ;
  assign n30584 = n30582 ^ n28818 ;
  assign n30583 = n30582 ^ n30574 ;
  assign n30585 = n30584 ^ n30583 ;
  assign n30586 = n30579 & ~n30585 ;
  assign n30587 = n30586 ^ n30584 ;
  assign n30653 = n30587 ^ n29575 ;
  assign n30835 = n30653 ^ x94 ;
  assign n30796 = n30795 ^ n30654 ;
  assign n30797 = ~n30655 & n30796 ;
  assign n30798 = n30797 ^ x95 ;
  assign n30836 = n30835 ^ n30798 ;
  assign n30908 = n30892 ^ n30836 ;
  assign n30909 = n30908 ^ n30540 ;
  assign n31262 = n30991 ^ n30909 ;
  assign n31263 = n29967 & n31262 ;
  assign n31264 = n31263 ^ n30540 ;
  assign n31265 = n31264 ^ n29239 ;
  assign n31269 = n31268 ^ n31265 ;
  assign n31271 = n31269 ^ x8 ;
  assign n31270 = n31269 ^ n31254 ;
  assign n31272 = n31271 ^ n31270 ;
  assign n31273 = ~n31259 & n31272 ;
  assign n31274 = n31273 ^ n31271 ;
  assign n31275 = n31274 ^ x23 ;
  assign n31276 = ~n31261 & n31275 ;
  assign n31287 = n31269 ^ x23 ;
  assign n31288 = n31274 & ~n31287 ;
  assign n31289 = n31288 ^ x23 ;
  assign n31290 = n31289 ^ x22 ;
  assign n30893 = n30836 & n30892 ;
  assign n30799 = n30798 ^ n30653 ;
  assign n30800 = n30798 ^ x94 ;
  assign n30801 = ~n30799 & n30800 ;
  assign n30802 = n30801 ^ x94 ;
  assign n30833 = n30802 ^ x93 ;
  assign n30421 = n30420 ^ n30411 ;
  assign n30422 = ~n30412 & n30421 ;
  assign n30423 = n30422 ^ n30013 ;
  assign n30409 = n30234 ^ n30232 ;
  assign n30408 = n29855 ^ n29638 ;
  assign n30410 = n30409 ^ n30408 ;
  assign n30424 = n30423 ^ n30410 ;
  assign n30425 = n30424 ^ n29855 ;
  assign n30589 = n30425 ^ n29575 ;
  assign n30588 = n30582 ^ n30425 ;
  assign n30590 = n30589 ^ n30588 ;
  assign n30591 = n30587 & n30590 ;
  assign n30592 = n30591 ^ n30589 ;
  assign n30803 = n30592 ^ n29618 ;
  assign n30834 = n30833 ^ n30803 ;
  assign n30995 = n30893 ^ n30834 ;
  assign n31281 = n30995 ^ n30440 ;
  assign n30992 = n30991 ^ n30908 ;
  assign n30993 = n30909 & n30992 ;
  assign n30994 = n30993 ^ n30540 ;
  assign n31282 = n31281 ^ n30994 ;
  assign n31283 = ~n29811 & ~n31282 ;
  assign n31284 = n31283 ^ n30440 ;
  assign n31285 = n31284 ^ n29246 ;
  assign n31277 = n31268 ^ n31264 ;
  assign n31278 = n31268 ^ n29239 ;
  assign n31279 = ~n31277 & n31278 ;
  assign n31280 = n31279 ^ n29239 ;
  assign n31286 = n31285 ^ n31280 ;
  assign n31291 = n31290 ^ n31286 ;
  assign n31292 = ~n31276 & ~n31291 ;
  assign n31302 = n31289 ^ n31286 ;
  assign n31303 = n31290 & n31302 ;
  assign n31304 = n31303 ^ x22 ;
  assign n31296 = n31284 ^ n31280 ;
  assign n31297 = n31285 & ~n31296 ;
  assign n31298 = n31297 ^ n29246 ;
  assign n31299 = n31298 ^ n29145 ;
  assign n30996 = n30995 ^ n30994 ;
  assign n30894 = n30834 & ~n30893 ;
  assign n30804 = n30803 ^ n30802 ;
  assign n30599 = n30236 ^ n30235 ;
  assign n30600 = n30599 ^ n30030 ;
  assign n30596 = n30423 ^ n30409 ;
  assign n30597 = ~n30410 & ~n30596 ;
  assign n30598 = n30597 ^ n30423 ;
  assign n30601 = n30600 ^ n30598 ;
  assign n30602 = n30601 ^ n30031 ;
  assign n30426 = n30425 ^ n29618 ;
  assign n30593 = n30426 & n30592 ;
  assign n30594 = n30593 ^ n29618 ;
  assign n30595 = n30594 ^ n28839 ;
  assign n30651 = n30602 ^ n30595 ;
  assign n30805 = n30651 ^ x93 ;
  assign n30806 = n30805 ^ n30651 ;
  assign n30807 = n30806 ^ n30802 ;
  assign n30808 = n30804 & n30807 ;
  assign n30809 = n30808 ^ n30805 ;
  assign n30832 = n30809 ^ x92 ;
  assign n30906 = n30894 ^ n30832 ;
  assign n30997 = n30906 ^ n30440 ;
  assign n30998 = n30997 ^ n30994 ;
  assign n30999 = n30998 ^ n30906 ;
  assign n31000 = ~n30996 & n30999 ;
  assign n31001 = n31000 ^ n30997 ;
  assign n31293 = n31001 ^ n30552 ;
  assign n31294 = ~n29891 & ~n31293 ;
  assign n31295 = n31294 ^ n30552 ;
  assign n31300 = n31299 ^ n31295 ;
  assign n31301 = n31300 ^ x21 ;
  assign n31305 = n31304 ^ n31301 ;
  assign n31306 = n31292 & ~n31305 ;
  assign n31316 = n31298 ^ n31295 ;
  assign n31317 = ~n31299 & n31316 ;
  assign n31318 = n31317 ^ n29145 ;
  assign n30895 = n30832 & ~n30894 ;
  assign n30603 = n30602 ^ n30594 ;
  assign n30604 = ~n30595 & n30603 ;
  assign n30605 = n30604 ^ n28839 ;
  assign n30813 = n30605 ^ n29632 ;
  assign n30608 = n30599 ^ n30598 ;
  assign n30609 = ~n30600 & ~n30608 ;
  assign n30610 = n30609 ^ n30030 ;
  assign n30606 = n30238 ^ n30237 ;
  assign n30607 = n30606 ^ n29876 ;
  assign n30611 = n30610 ^ n30607 ;
  assign n30612 = n30611 ^ n29877 ;
  assign n30814 = n30813 ^ n30612 ;
  assign n30652 = n30651 ^ x92 ;
  assign n30810 = n30652 & ~n30809 ;
  assign n30811 = n30810 ^ x92 ;
  assign n30812 = n30811 ^ x91 ;
  assign n30831 = n30814 ^ n30812 ;
  assign n30905 = n30895 ^ n30831 ;
  assign n31311 = n30905 ^ n30438 ;
  assign n30907 = n30906 ^ n30552 ;
  assign n31002 = n30907 & n31001 ;
  assign n31003 = n31002 ^ n30552 ;
  assign n31312 = n31311 ^ n31003 ;
  assign n31313 = n29806 & ~n31312 ;
  assign n31314 = n31313 ^ n30438 ;
  assign n31315 = n31314 ^ n29269 ;
  assign n31319 = n31318 ^ n31315 ;
  assign n31320 = n31319 ^ x20 ;
  assign n31307 = n31304 ^ n31300 ;
  assign n31308 = n31304 ^ x21 ;
  assign n31309 = n31307 & n31308 ;
  assign n31310 = n31309 ^ x21 ;
  assign n31321 = n31320 ^ n31310 ;
  assign n31322 = ~n31306 & ~n31321 ;
  assign n31333 = n31319 ^ n31310 ;
  assign n31334 = n31320 & ~n31333 ;
  assign n31335 = n31334 ^ x20 ;
  assign n31336 = n31335 ^ x19 ;
  assign n31327 = n31318 ^ n31314 ;
  assign n31328 = n31318 ^ n29269 ;
  assign n31329 = ~n31327 & n31328 ;
  assign n31330 = n31329 ^ n29269 ;
  assign n31331 = n31330 ^ n29282 ;
  assign n30896 = n30831 & n30895 ;
  assign n30613 = n30612 ^ n30605 ;
  assign n30614 = n30612 ^ n29632 ;
  assign n30615 = n30613 & ~n30614 ;
  assign n30616 = n30615 ^ n29632 ;
  assign n30818 = n30616 ^ n28854 ;
  assign n30622 = n30240 ^ n30239 ;
  assign n30621 = n29868 ^ n29685 ;
  assign n30623 = n30622 ^ n30621 ;
  assign n30617 = n30610 ^ n30606 ;
  assign n30618 = n30610 ^ n29876 ;
  assign n30619 = n30617 & ~n30618 ;
  assign n30620 = n30619 ^ n29876 ;
  assign n30624 = n30623 ^ n30620 ;
  assign n30625 = n30624 ^ n29868 ;
  assign n30819 = n30818 ^ n30625 ;
  assign n30829 = n30819 ^ x90 ;
  assign n30815 = n30814 ^ n30811 ;
  assign n30816 = n30812 & ~n30815 ;
  assign n30817 = n30816 ^ x91 ;
  assign n30830 = n30829 ^ n30817 ;
  assign n31008 = n30896 ^ n30830 ;
  assign n31323 = n31008 ^ n30435 ;
  assign n31004 = n31003 ^ n30905 ;
  assign n31005 = n31003 ^ n30438 ;
  assign n31006 = n31004 & n31005 ;
  assign n31007 = n31006 ^ n30438 ;
  assign n31324 = n31323 ^ n31007 ;
  assign n31325 = ~n29884 & ~n31324 ;
  assign n31326 = n31325 ^ n30435 ;
  assign n31332 = n31331 ^ n31326 ;
  assign n31337 = n31336 ^ n31332 ;
  assign n31338 = ~n31322 & ~n31337 ;
  assign n31348 = n31335 ^ n31332 ;
  assign n31349 = n31336 & n31348 ;
  assign n31350 = n31349 ^ x19 ;
  assign n31351 = n31350 ^ x18 ;
  assign n31343 = n31326 ^ n29282 ;
  assign n31344 = n31330 ^ n31326 ;
  assign n31345 = ~n31343 & n31344 ;
  assign n31346 = n31345 ^ n29282 ;
  assign n31009 = n31008 ^ n31007 ;
  assign n30820 = n30819 ^ n30817 ;
  assign n30626 = n30625 ^ n30616 ;
  assign n30627 = n30625 ^ n28854 ;
  assign n30628 = ~n30626 & n30627 ;
  assign n30629 = n30628 ^ n28854 ;
  assign n30821 = n30629 ^ n29703 ;
  assign n30634 = n30243 ^ n30241 ;
  assign n30633 = n30194 ^ n29870 ;
  assign n30635 = n30634 ^ n30633 ;
  assign n30630 = n30621 ^ n30620 ;
  assign n30631 = ~n30623 & n30630 ;
  assign n30632 = n30631 ^ n30622 ;
  assign n30636 = n30635 ^ n30632 ;
  assign n30637 = n30636 ^ n29871 ;
  assign n30822 = n30821 ^ n30637 ;
  assign n30823 = n30822 ^ x90 ;
  assign n30824 = n30823 ^ n30817 ;
  assign n30825 = n30824 ^ n30822 ;
  assign n30826 = n30820 & n30825 ;
  assign n30827 = n30826 ^ n30823 ;
  assign n31010 = n30827 ^ x89 ;
  assign n30897 = ~n30830 & n30896 ;
  assign n31011 = n31010 ^ n30897 ;
  assign n31012 = n31011 ^ n30435 ;
  assign n31013 = n31012 ^ n31011 ;
  assign n31014 = n31013 ^ n31007 ;
  assign n31015 = ~n31009 & ~n31014 ;
  assign n31016 = n31015 ^ n31012 ;
  assign n31339 = n31016 ^ n30432 ;
  assign n31340 = ~n30388 & n31339 ;
  assign n31341 = n31340 ^ n30432 ;
  assign n31342 = n31341 ^ n29293 ;
  assign n31347 = n31346 ^ n31342 ;
  assign n31352 = n31351 ^ n31347 ;
  assign n31353 = ~n31338 & ~n31352 ;
  assign n31364 = n31350 ^ n31347 ;
  assign n31365 = n31351 & ~n31364 ;
  assign n31366 = n31365 ^ x18 ;
  assign n31357 = n31346 ^ n31341 ;
  assign n31358 = n31346 ^ n29293 ;
  assign n31359 = n31357 & ~n31358 ;
  assign n31360 = n31359 ^ n29293 ;
  assign n31361 = n31360 ^ n29430 ;
  assign n30898 = n30897 ^ n30822 ;
  assign n30901 = ~n30827 & ~n30898 ;
  assign n30828 = n30827 ^ n30822 ;
  assign n30899 = n30898 ^ n30828 ;
  assign n30900 = x89 & ~n30899 ;
  assign n30902 = n30901 ^ n30900 ;
  assign n30647 = n30198 ^ n29703 ;
  assign n30643 = n30245 ^ n30244 ;
  assign n30644 = n30643 ^ n30196 ;
  assign n30645 = n30644 ^ n30634 ;
  assign n30641 = n30633 ^ n30632 ;
  assign n30642 = n30635 & ~n30641 ;
  assign n30646 = n30645 ^ n30642 ;
  assign n30648 = n30647 ^ n30646 ;
  assign n30649 = n30648 ^ x88 ;
  assign n30638 = n30637 ^ n30629 ;
  assign n30639 = n30637 ^ n29703 ;
  assign n30640 = n30638 & ~n30639 ;
  assign n30650 = n30649 ^ n30640 ;
  assign n30903 = n30902 ^ n30650 ;
  assign n31018 = n30903 ^ n30432 ;
  assign n31017 = n31011 ^ n30903 ;
  assign n31019 = n31018 ^ n31017 ;
  assign n31020 = n31016 & ~n31019 ;
  assign n31021 = n31020 ^ n31018 ;
  assign n31354 = n31021 ^ n30428 ;
  assign n31355 = n30390 & n31354 ;
  assign n31356 = n31355 ^ n30428 ;
  assign n31362 = n31361 ^ n31356 ;
  assign n31363 = n31362 ^ x17 ;
  assign n31367 = n31366 ^ n31363 ;
  assign n31368 = ~n31353 & ~n31367 ;
  assign n31377 = n31366 ^ n31362 ;
  assign n31378 = n31366 ^ x17 ;
  assign n31379 = n31377 & n31378 ;
  assign n31380 = n31379 ^ x17 ;
  assign n31381 = n31380 ^ x16 ;
  assign n31372 = n31356 ^ n29430 ;
  assign n31373 = n31360 ^ n31356 ;
  assign n31374 = n31372 & n31373 ;
  assign n31375 = n31374 ^ n29430 ;
  assign n30904 = n30903 ^ n30428 ;
  assign n31022 = ~n30904 & ~n31021 ;
  assign n31023 = n31022 ^ n30428 ;
  assign n30407 = n30406 ^ n30404 ;
  assign n31024 = n31023 ^ n30407 ;
  assign n31369 = n30000 & n31024 ;
  assign n31370 = n31369 ^ n30404 ;
  assign n31371 = n31370 ^ n29495 ;
  assign n31376 = n31375 ^ n31371 ;
  assign n31382 = n31381 ^ n31376 ;
  assign n31383 = n31368 & ~n31382 ;
  assign n31384 = n31380 ^ n31376 ;
  assign n31402 = n31381 & n31384 ;
  assign n31393 = n31375 ^ n31370 ;
  assign n31394 = n31375 ^ n29495 ;
  assign n31395 = n31393 & n31394 ;
  assign n31396 = n31395 ^ n29495 ;
  assign n31397 = n31396 ^ n29528 ;
  assign n31388 = n30859 ^ n30406 ;
  assign n31389 = n31388 ^ n30573 ;
  assign n31385 = n31023 ^ n30404 ;
  assign n31386 = n30407 & n31385 ;
  assign n31387 = n31386 ^ n30406 ;
  assign n31390 = n31389 ^ n31387 ;
  assign n31391 = n30004 & n31390 ;
  assign n31392 = n31391 ^ n30573 ;
  assign n31398 = n31397 ^ n31392 ;
  assign n31399 = n31398 ^ x16 ;
  assign n31403 = n31402 ^ n31399 ;
  assign n31404 = n31403 ^ x31 ;
  assign n31405 = n31383 & n31404 ;
  assign n31423 = n31398 ^ x31 ;
  assign n31424 = ~n31403 & n31423 ;
  assign n31425 = n31424 ^ x31 ;
  assign n31417 = n31392 ^ n29528 ;
  assign n31418 = n31396 ^ n31392 ;
  assign n31419 = n31417 & n31418 ;
  assign n31420 = n31419 ^ n29528 ;
  assign n31412 = n30862 ^ n30860 ;
  assign n31406 = n31388 ^ n31387 ;
  assign n31407 = n30580 ^ n30573 ;
  assign n31408 = n31407 ^ n30580 ;
  assign n31409 = n31408 ^ n31387 ;
  assign n31410 = n31406 & n31409 ;
  assign n31411 = n31410 ^ n31407 ;
  assign n31413 = n31412 ^ n31411 ;
  assign n31414 = n30013 & n31413 ;
  assign n31415 = n31414 ^ n30580 ;
  assign n31416 = n31415 ^ n29576 ;
  assign n31421 = n31420 ^ n31416 ;
  assign n31422 = n31421 ^ x30 ;
  assign n31426 = n31425 ^ n31422 ;
  assign n31427 = n31405 & ~n31426 ;
  assign n31439 = n31412 ^ n30580 ;
  assign n31440 = ~n31411 & ~n31439 ;
  assign n31441 = n31440 ^ n30580 ;
  assign n31437 = n30864 ^ n30863 ;
  assign n31438 = n31437 ^ n30424 ;
  assign n31442 = n31441 ^ n31438 ;
  assign n31443 = ~n30408 & ~n31442 ;
  assign n31444 = n31443 ^ n30424 ;
  assign n31432 = n31420 ^ n31415 ;
  assign n31433 = n31420 ^ n29576 ;
  assign n31434 = n31432 & ~n31433 ;
  assign n31435 = n31434 ^ n29576 ;
  assign n31436 = n31435 ^ n29638 ;
  assign n31445 = n31444 ^ n31436 ;
  assign n31446 = n31445 ^ x29 ;
  assign n31428 = n31425 ^ n31421 ;
  assign n31429 = n31425 ^ x30 ;
  assign n31430 = n31428 & n31429 ;
  assign n31431 = n31430 ^ x30 ;
  assign n31447 = n31446 ^ n31431 ;
  assign n31448 = ~n31427 & ~n31447 ;
  assign n31466 = n31445 ^ n31431 ;
  assign n31467 = n31446 & ~n31466 ;
  assign n31468 = n31467 ^ x29 ;
  assign n31449 = n31444 ^ n31435 ;
  assign n31454 = n30866 ^ n30865 ;
  assign n31455 = n31454 ^ n30601 ;
  assign n31450 = n31441 ^ n31437 ;
  assign n31451 = n31441 ^ n30424 ;
  assign n31452 = ~n31450 & ~n31451 ;
  assign n31453 = n31452 ^ n30424 ;
  assign n31456 = n31455 ^ n31453 ;
  assign n31457 = ~n30030 & ~n31456 ;
  assign n31458 = n31457 ^ n30601 ;
  assign n31459 = n31458 ^ n29638 ;
  assign n31460 = n31459 ^ n31458 ;
  assign n31461 = n31460 ^ n31435 ;
  assign n31462 = n31449 & ~n31461 ;
  assign n31463 = n31462 ^ n31459 ;
  assign n31464 = n31463 ^ n29649 ;
  assign n31465 = n31464 ^ x28 ;
  assign n31469 = n31468 ^ n31465 ;
  assign n31470 = ~n31448 & n31469 ;
  assign n31471 = n31468 ^ n31464 ;
  assign n31489 = n31468 ^ x28 ;
  assign n31490 = ~n31471 & n31489 ;
  assign n31482 = n30868 ^ n30867 ;
  assign n31476 = n31454 ^ n31453 ;
  assign n31477 = n30611 ^ n30601 ;
  assign n31478 = n31477 ^ n30611 ;
  assign n31479 = n31478 ^ n31453 ;
  assign n31480 = n31476 & ~n31479 ;
  assign n31481 = n31480 ^ n31477 ;
  assign n31483 = n31482 ^ n31481 ;
  assign n31484 = n29876 & n31483 ;
  assign n31485 = n31484 ^ n30611 ;
  assign n31472 = n31458 ^ n29649 ;
  assign n31473 = n31463 & ~n31472 ;
  assign n31474 = n31473 ^ n29649 ;
  assign n31475 = n31474 ^ n29635 ;
  assign n31486 = n31485 ^ n31475 ;
  assign n31487 = n31486 ^ x28 ;
  assign n31491 = n31490 ^ n31487 ;
  assign n31492 = n31491 ^ x27 ;
  assign n31493 = ~n31470 & ~n31492 ;
  assign n31507 = n31485 ^ n29635 ;
  assign n31508 = n31485 ^ n31474 ;
  assign n31509 = ~n31507 & n31508 ;
  assign n31510 = n31509 ^ n29635 ;
  assign n31502 = n30871 ^ n30869 ;
  assign n31498 = n30624 ^ n30611 ;
  assign n31497 = n31482 ^ n30624 ;
  assign n31499 = n31498 ^ n31497 ;
  assign n31500 = n31481 & n31499 ;
  assign n31501 = n31500 ^ n31498 ;
  assign n31503 = n31502 ^ n31501 ;
  assign n31504 = ~n30621 & ~n31503 ;
  assign n31505 = n31504 ^ n30624 ;
  assign n31506 = n31505 ^ n29685 ;
  assign n31511 = n31510 ^ n31506 ;
  assign n31512 = n31511 ^ x26 ;
  assign n31494 = n31486 ^ x27 ;
  assign n31495 = ~n31491 & n31494 ;
  assign n31496 = n31495 ^ x27 ;
  assign n31513 = n31512 ^ n31496 ;
  assign n31514 = n31493 & ~n31513 ;
  assign n31530 = n31511 ^ n31496 ;
  assign n31531 = n31512 & ~n31530 ;
  assign n31532 = n31531 ^ x26 ;
  assign n31522 = n31502 ^ n30624 ;
  assign n31523 = n31501 & ~n31522 ;
  assign n31524 = n31523 ^ n30624 ;
  assign n31520 = n30873 ^ n30872 ;
  assign n31521 = n31520 ^ n30636 ;
  assign n31525 = n31524 ^ n31521 ;
  assign n31526 = n30633 & n31525 ;
  assign n31527 = n31526 ^ n30636 ;
  assign n31515 = n31510 ^ n31505 ;
  assign n31516 = n31510 ^ n29685 ;
  assign n31517 = n31515 & n31516 ;
  assign n31518 = n31517 ^ n29685 ;
  assign n31519 = n31518 ^ n29709 ;
  assign n31528 = n31527 ^ n31519 ;
  assign n31529 = n31528 ^ x25 ;
  assign n31533 = n31532 ^ n31529 ;
  assign n31576 = n31514 & ~n31533 ;
  assign n31568 = n30875 ^ n30646 ;
  assign n31569 = n31568 ^ n30874 ;
  assign n31570 = n31569 ^ n31520 ;
  assign n31565 = n31524 ^ n31520 ;
  assign n31566 = n31524 ^ n30636 ;
  assign n31567 = ~n31565 & n31566 ;
  assign n31571 = n31570 ^ n31567 ;
  assign n31572 = ~n30196 & ~n31571 ;
  assign n31562 = n29751 ^ n29709 ;
  assign n31563 = n31562 ^ n30646 ;
  assign n31564 = n31563 ^ n610 ;
  assign n31573 = n31572 ^ n31564 ;
  assign n31559 = n31527 ^ n31518 ;
  assign n31560 = n31527 ^ n29709 ;
  assign n31561 = ~n31559 & ~n31560 ;
  assign n31574 = n31573 ^ n31561 ;
  assign n31556 = n31532 ^ n31528 ;
  assign n31557 = n31532 ^ x25 ;
  assign n31558 = ~n31556 & n31557 ;
  assign n31575 = n31574 ^ n31558 ;
  assign n31577 = n31576 ^ n31575 ;
  assign n31534 = n31533 ^ n31514 ;
  assign n31535 = n31534 ^ n31071 ;
  assign n31536 = n31513 ^ n31493 ;
  assign n31537 = n31536 ^ n31060 ;
  assign n31538 = n31447 ^ n31427 ;
  assign n31539 = ~n31026 & ~n31538 ;
  assign n31540 = n31539 ^ n31034 ;
  assign n31541 = n31469 ^ n31448 ;
  assign n31542 = n31541 ^ n31539 ;
  assign n31543 = ~n31540 & n31542 ;
  assign n31544 = n31543 ^ n31034 ;
  assign n31545 = n31544 ^ n31049 ;
  assign n31546 = n31492 ^ n31470 ;
  assign n31547 = n31546 ^ n31544 ;
  assign n31548 = n31545 & ~n31547 ;
  assign n31549 = n31548 ^ n31049 ;
  assign n31550 = n31549 ^ n31536 ;
  assign n31551 = ~n31537 & n31550 ;
  assign n31552 = n31551 ^ n31060 ;
  assign n31553 = n31552 ^ n31534 ;
  assign n31554 = ~n31535 & n31553 ;
  assign n31555 = n31554 ^ n31071 ;
  assign n31578 = n31577 ^ n31555 ;
  assign n31609 = n31555 ^ n31088 ;
  assign n31582 = ~n31578 & ~n31609 ;
  assign n31579 = n31088 ^ n31029 ;
  assign n31583 = n31582 ^ n31579 ;
  assign n31584 = n31031 & n31583 ;
  assign n31585 = n31584 ^ n31030 ;
  assign n31587 = n31586 ^ n31585 ;
  assign n31588 = n31136 ^ n31118 ;
  assign n31589 = n31588 ^ n31136 ;
  assign n31590 = n31589 ^ n31585 ;
  assign n31591 = n31587 & n31590 ;
  assign n31592 = n31591 ^ n31588 ;
  assign n31602 = n31592 ^ n31053 ;
  assign n31603 = n30457 & ~n31602 ;
  assign n31604 = n31603 ^ n31136 ;
  assign n31605 = n31604 ^ n30287 ;
  assign n31653 = n31586 ^ n31118 ;
  assign n31654 = n31653 ^ n31585 ;
  assign n31655 = n30460 & ~n31654 ;
  assign n31656 = n31655 ^ n31118 ;
  assign n31610 = n31609 ^ n31577 ;
  assign n31611 = ~n30465 & ~n31610 ;
  assign n31612 = n31611 ^ n31088 ;
  assign n31613 = n31612 ^ n30301 ;
  assign n31614 = n31552 ^ n31535 ;
  assign n31615 = ~n30468 & ~n31614 ;
  assign n31616 = n31615 ^ n31071 ;
  assign n31617 = n31616 ^ n30305 ;
  assign n31618 = n31549 ^ n31537 ;
  assign n31619 = ~n30471 & ~n31618 ;
  assign n31620 = n31619 ^ n31060 ;
  assign n31621 = n31620 ^ n30308 ;
  assign n31628 = n31538 ^ n31026 ;
  assign n31629 = n30925 & ~n31628 ;
  assign n31630 = n31629 ^ n31026 ;
  assign n31631 = ~n30318 & n31630 ;
  assign n31625 = n31541 ^ n31540 ;
  assign n31626 = n30479 & ~n31625 ;
  assign n31627 = n31626 ^ n31034 ;
  assign n31632 = n31631 ^ n31627 ;
  assign n31633 = n31631 ^ n30321 ;
  assign n31634 = ~n31632 & ~n31633 ;
  assign n31635 = n31634 ^ n30321 ;
  assign n31622 = n31546 ^ n31545 ;
  assign n31623 = ~n30474 & n31622 ;
  assign n31624 = n31623 ^ n31049 ;
  assign n31636 = n31635 ^ n31624 ;
  assign n31637 = n31635 ^ n30314 ;
  assign n31638 = n31636 & ~n31637 ;
  assign n31639 = n31638 ^ n30314 ;
  assign n31640 = n31639 ^ n31620 ;
  assign n31641 = n31621 & ~n31640 ;
  assign n31642 = n31641 ^ n30308 ;
  assign n31643 = n31642 ^ n31616 ;
  assign n31644 = ~n31617 & ~n31643 ;
  assign n31645 = n31644 ^ n30305 ;
  assign n31646 = n31645 ^ n31612 ;
  assign n31647 = n31613 & ~n31646 ;
  assign n31648 = n31647 ^ n30301 ;
  assign n31606 = n31583 ^ n31030 ;
  assign n31607 = ~n30462 & ~n31606 ;
  assign n31608 = n31607 ^ n31030 ;
  assign n31649 = n31648 ^ n31608 ;
  assign n31650 = n31648 ^ n30297 ;
  assign n31651 = n31649 & ~n31650 ;
  assign n31652 = n31651 ^ n30297 ;
  assign n31657 = n31656 ^ n31652 ;
  assign n31685 = n31652 ^ n30292 ;
  assign n31661 = ~n31657 & n31685 ;
  assign n31658 = n31604 ^ n30292 ;
  assign n31662 = n31661 ^ n31658 ;
  assign n31663 = n31605 & n31662 ;
  assign n31664 = n31663 ^ n30287 ;
  assign n31681 = n31664 ^ n30285 ;
  assign n31593 = n31069 ^ n31053 ;
  assign n31594 = n31593 ^ n31136 ;
  assign n31596 = n31594 ^ n31069 ;
  assign n31597 = n31592 & ~n31596 ;
  assign n31598 = n31597 ^ n31069 ;
  assign n31599 = n31598 ^ n31151 ;
  assign n31600 = ~n30510 & n31599 ;
  assign n31601 = n31600 ^ n31151 ;
  assign n31682 = n31681 ^ n31601 ;
  assign n31683 = n31682 ^ x238 ;
  assign n31686 = n31685 ^ n31656 ;
  assign n31687 = n31686 ^ x224 ;
  assign n31690 = n31645 ^ n31613 ;
  assign n31691 = n31690 ^ x226 ;
  assign n31705 = n31639 ^ n30308 ;
  assign n31706 = n31705 ^ n31620 ;
  assign n31700 = n31637 ^ n31624 ;
  assign n31693 = n30926 ^ n30317 ;
  assign n31694 = n31693 ^ n31629 ;
  assign n31695 = x231 & ~n31694 ;
  assign n31692 = n31633 ^ n31627 ;
  assign n31696 = n31695 ^ n31692 ;
  assign n31697 = n31695 ^ x230 ;
  assign n31698 = n31696 & n31697 ;
  assign n31699 = n31698 ^ x230 ;
  assign n31701 = n31700 ^ n31699 ;
  assign n31702 = n31700 ^ x229 ;
  assign n31703 = n31701 & ~n31702 ;
  assign n31704 = n31703 ^ x229 ;
  assign n31707 = n31706 ^ n31704 ;
  assign n31708 = n31642 ^ n31617 ;
  assign n31709 = n31708 ^ x228 ;
  assign n31710 = n31709 ^ n31708 ;
  assign n31711 = n31710 ^ n31704 ;
  assign n31712 = ~n31707 & n31711 ;
  assign n31713 = n31712 ^ n31709 ;
  assign n31715 = n31690 ^ x227 ;
  assign n31714 = n31708 ^ n31690 ;
  assign n31716 = n31715 ^ n31714 ;
  assign n31717 = n31713 & ~n31716 ;
  assign n31718 = n31717 ^ n31715 ;
  assign n31719 = ~n31691 & n31718 ;
  assign n31720 = n31719 ^ x226 ;
  assign n31688 = n31608 ^ n30297 ;
  assign n31689 = n31688 ^ n31648 ;
  assign n31721 = n31720 ^ n31689 ;
  assign n31722 = n31686 ^ x225 ;
  assign n31723 = n31722 ^ n31686 ;
  assign n31724 = n31723 ^ n31689 ;
  assign n31725 = n31721 & ~n31724 ;
  assign n31726 = n31725 ^ n31722 ;
  assign n31727 = n31687 & ~n31726 ;
  assign n31728 = n31727 ^ x224 ;
  assign n31684 = n31662 ^ n30287 ;
  assign n31729 = n31728 ^ n31684 ;
  assign n31730 = n31728 ^ x239 ;
  assign n31731 = ~n31729 & n31730 ;
  assign n31732 = n31731 ^ x239 ;
  assign n31733 = n31732 ^ n31682 ;
  assign n31734 = n31683 & ~n31733 ;
  assign n31735 = n31734 ^ x238 ;
  assign n31665 = n31664 ^ n31601 ;
  assign n31677 = n31601 ^ n30285 ;
  assign n31678 = ~n31665 & ~n31677 ;
  assign n31666 = n31085 ^ n31070 ;
  assign n31668 = n31666 ^ n31151 ;
  assign n31667 = n31666 ^ n31593 ;
  assign n31669 = n31668 ^ n31667 ;
  assign n31670 = n31598 & n31669 ;
  assign n31671 = n31670 ^ n31668 ;
  assign n31672 = n31671 ^ n31165 ;
  assign n31673 = ~n30455 & n31672 ;
  assign n31674 = n31673 ^ n31165 ;
  assign n31675 = n31674 ^ n30285 ;
  assign n31679 = n31678 ^ n31675 ;
  assign n31680 = n31679 ^ n30279 ;
  assign n31736 = n31735 ^ n31680 ;
  assign n31743 = n31101 ^ n31086 ;
  assign n31744 = n31743 ^ n31185 ;
  assign n31740 = n31666 ^ n31165 ;
  assign n31741 = n31671 & ~n31740 ;
  assign n31742 = n31741 ^ n31165 ;
  assign n31745 = n31744 ^ n31742 ;
  assign n31746 = ~n30452 & ~n31745 ;
  assign n31747 = n31746 ^ n31185 ;
  assign n31748 = n31747 ^ n30275 ;
  assign n31737 = n31674 ^ n30279 ;
  assign n31738 = n31679 & n31737 ;
  assign n31739 = n31738 ^ n30279 ;
  assign n31749 = n31748 ^ n31739 ;
  assign n31750 = n31749 ^ x237 ;
  assign n31751 = n31750 ^ n31680 ;
  assign n31752 = n31751 ^ n31749 ;
  assign n31753 = ~n31736 & n31752 ;
  assign n31754 = n31753 ^ n31750 ;
  assign n31765 = n31115 ^ n31102 ;
  assign n31759 = n31743 ^ n31742 ;
  assign n31760 = n31200 ^ n31185 ;
  assign n31761 = n31760 ^ n31200 ;
  assign n31762 = n31761 ^ n31742 ;
  assign n31763 = n31759 & ~n31762 ;
  assign n31764 = n31763 ^ n31760 ;
  assign n31766 = n31765 ^ n31764 ;
  assign n31767 = n30450 & ~n31766 ;
  assign n31768 = n31767 ^ n31200 ;
  assign n31755 = n31747 ^ n31739 ;
  assign n31756 = n31748 & n31755 ;
  assign n31757 = n31756 ^ n30275 ;
  assign n31758 = n31757 ^ n29950 ;
  assign n31769 = n31768 ^ n31758 ;
  assign n31771 = n31769 ^ x236 ;
  assign n31770 = n31769 ^ n31749 ;
  assign n31772 = n31771 ^ n31770 ;
  assign n31773 = n31754 & ~n31772 ;
  assign n31774 = n31773 ^ n31771 ;
  assign n32097 = n31769 ^ x235 ;
  assign n32098 = n31774 & ~n32097 ;
  assign n32099 = n32098 ^ x235 ;
  assign n32100 = n32099 ^ x234 ;
  assign n31969 = n31768 ^ n31757 ;
  assign n31821 = n31132 ^ n31116 ;
  assign n31964 = n31821 ^ n31217 ;
  assign n31822 = n31765 ^ n31200 ;
  assign n31823 = ~n31764 & ~n31822 ;
  assign n31824 = n31823 ^ n31200 ;
  assign n31965 = n31964 ^ n31824 ;
  assign n31966 = n30446 & ~n31965 ;
  assign n31967 = n31966 ^ n31217 ;
  assign n31970 = n31967 ^ n29950 ;
  assign n31971 = n31970 ^ n31967 ;
  assign n31972 = n31971 ^ n31768 ;
  assign n31973 = n31969 & ~n31972 ;
  assign n31974 = n31973 ^ n31970 ;
  assign n32101 = n31974 ^ n29904 ;
  assign n32102 = n32101 ^ n32099 ;
  assign n32103 = n32100 & ~n32102 ;
  assign n32104 = n32103 ^ x234 ;
  assign n32196 = n32104 ^ x233 ;
  assign n31968 = n31967 ^ n29904 ;
  assign n31975 = n31968 & n31974 ;
  assign n31976 = n31975 ^ n29904 ;
  assign n31825 = n31824 ^ n31821 ;
  assign n31826 = n31232 ^ n31217 ;
  assign n31827 = n31826 ^ n31232 ;
  assign n31828 = n31827 ^ n31821 ;
  assign n31829 = ~n31825 & n31828 ;
  assign n31830 = n31829 ^ n31826 ;
  assign n31819 = n31149 ^ n31133 ;
  assign n31876 = n31830 ^ n31819 ;
  assign n31961 = n30444 & n31876 ;
  assign n31962 = n31961 ^ n31232 ;
  assign n31963 = n31962 ^ n29900 ;
  assign n32095 = n31976 ^ n31963 ;
  assign n32197 = n32196 ^ n32095 ;
  assign n31775 = n31774 ^ x235 ;
  assign n31776 = n31713 ^ x227 ;
  assign n31777 = n31694 ^ x231 ;
  assign n31778 = n31692 ^ x230 ;
  assign n31779 = n31778 ^ n31695 ;
  assign n31780 = n31777 & n31779 ;
  assign n31781 = n31699 ^ x229 ;
  assign n31782 = n31781 ^ n31700 ;
  assign n31783 = n31780 & n31782 ;
  assign n31784 = n31706 ^ x228 ;
  assign n31785 = n31784 ^ n31704 ;
  assign n31786 = ~n31783 & n31785 ;
  assign n31787 = n31776 & ~n31786 ;
  assign n31788 = n31718 ^ x226 ;
  assign n31789 = ~n31787 & ~n31788 ;
  assign n31790 = n31689 ^ x225 ;
  assign n31791 = n31790 ^ n31720 ;
  assign n31792 = n31789 & ~n31791 ;
  assign n31793 = n31726 ^ x224 ;
  assign n31794 = ~n31792 & ~n31793 ;
  assign n31795 = n31684 ^ x239 ;
  assign n31796 = n31795 ^ n31728 ;
  assign n31797 = n31794 & ~n31796 ;
  assign n31798 = n31732 ^ n31683 ;
  assign n31799 = n31797 & ~n31798 ;
  assign n31800 = n31680 ^ x237 ;
  assign n31801 = n31800 ^ n31735 ;
  assign n31802 = n31799 & ~n31801 ;
  assign n31803 = n31754 ^ x236 ;
  assign n31804 = n31802 & n31803 ;
  assign n32192 = n31775 & n31804 ;
  assign n32193 = n32101 ^ x234 ;
  assign n32194 = n32193 ^ n32099 ;
  assign n32195 = n32192 & ~n32194 ;
  assign n32706 = n32197 ^ n32195 ;
  assign n31888 = n31305 ^ n31292 ;
  assign n31938 = n31888 ^ n31390 ;
  assign n31889 = n31291 ^ n31276 ;
  assign n31890 = n31889 ^ n31024 ;
  assign n31807 = n31260 ^ n31243 ;
  assign n31808 = n31807 ^ n31339 ;
  assign n31810 = n31227 ^ n31210 ;
  assign n31811 = n31810 ^ n31312 ;
  assign n31812 = n31209 ^ n31196 ;
  assign n31813 = n31812 ^ n31293 ;
  assign n31814 = n31195 ^ n31178 ;
  assign n31815 = n31814 ^ n31282 ;
  assign n31816 = n31177 ^ n31164 ;
  assign n31817 = n31816 ^ n31262 ;
  assign n31820 = n31819 ^ n31232 ;
  assign n31831 = ~n31820 & ~n31830 ;
  assign n31832 = n31831 ^ n31232 ;
  assign n31818 = n31163 ^ n31150 ;
  assign n31833 = n31832 ^ n31818 ;
  assign n31834 = n31816 ^ n31246 ;
  assign n31835 = n31834 ^ n31816 ;
  assign n31836 = n31835 ^ n31818 ;
  assign n31837 = ~n31833 & n31836 ;
  assign n31838 = n31837 ^ n31834 ;
  assign n31839 = ~n31817 & n31838 ;
  assign n31840 = n31839 ^ n31262 ;
  assign n31841 = n31840 ^ n31814 ;
  assign n31842 = n31815 & n31841 ;
  assign n31843 = n31842 ^ n31282 ;
  assign n31844 = n31843 ^ n31812 ;
  assign n31845 = n31813 & ~n31844 ;
  assign n31846 = n31845 ^ n31293 ;
  assign n31847 = n31846 ^ n31810 ;
  assign n31848 = n31811 & ~n31847 ;
  assign n31849 = n31848 ^ n31312 ;
  assign n31809 = n31242 ^ n31228 ;
  assign n31850 = n31849 ^ n31809 ;
  assign n31851 = n31339 ^ n31324 ;
  assign n31852 = n31851 ^ n31339 ;
  assign n31853 = n31852 ^ n31809 ;
  assign n31854 = n31850 & ~n31853 ;
  assign n31855 = n31854 ^ n31851 ;
  assign n31856 = ~n31808 & ~n31855 ;
  assign n31857 = n31856 ^ n31339 ;
  assign n31806 = n31275 ^ n31261 ;
  assign n31858 = n31857 ^ n31806 ;
  assign n31891 = n31889 ^ n31354 ;
  assign n31892 = n31891 ^ n31857 ;
  assign n31893 = n31892 ^ n31889 ;
  assign n31894 = n31858 & n31893 ;
  assign n31895 = n31894 ^ n31891 ;
  assign n31896 = ~n31890 & n31895 ;
  assign n31897 = n31896 ^ n31024 ;
  assign n31939 = n31938 ^ n31897 ;
  assign n32707 = n32706 ^ n31939 ;
  assign n32325 = n32194 ^ n32192 ;
  assign n31942 = n31895 ^ n31024 ;
  assign n32326 = n32325 ^ n31942 ;
  assign n31859 = n31858 ^ n31354 ;
  assign n31805 = n31804 ^ n31775 ;
  assign n31860 = n31859 ^ n31805 ;
  assign n31863 = n31809 ^ n31324 ;
  assign n31864 = n31863 ^ n31849 ;
  assign n31862 = n31801 ^ n31799 ;
  assign n31865 = n31864 ^ n31862 ;
  assign n31868 = n31798 ^ n31797 ;
  assign n31866 = n31846 ^ n31811 ;
  assign n31869 = n31868 ^ n31866 ;
  assign n31872 = n31838 ^ n31262 ;
  assign n31871 = n31791 ^ n31789 ;
  assign n31873 = n31872 ^ n31871 ;
  assign n31956 = n31818 ^ n31246 ;
  assign n31957 = n31956 ^ n31832 ;
  assign n32298 = n31957 ^ n31872 ;
  assign n31875 = n31786 ^ n31776 ;
  assign n31877 = n31876 ^ n31875 ;
  assign n31879 = n31782 ^ n31780 ;
  assign n31880 = n31879 ^ n31766 ;
  assign n32279 = n31779 ^ n31777 ;
  assign n31881 = n31777 ^ n31672 ;
  assign n31886 = n31321 ^ n31306 ;
  assign n31887 = n31886 ^ n31413 ;
  assign n31898 = n31897 ^ n31888 ;
  assign n31899 = n31413 ^ n31390 ;
  assign n31900 = n31899 ^ n31413 ;
  assign n31901 = n31900 ^ n31888 ;
  assign n31902 = ~n31898 & n31901 ;
  assign n31903 = n31902 ^ n31899 ;
  assign n31904 = n31887 & n31903 ;
  assign n31905 = n31904 ^ n31413 ;
  assign n31885 = n31337 ^ n31322 ;
  assign n31906 = n31905 ^ n31885 ;
  assign n31907 = n31456 ^ n31442 ;
  assign n31908 = n31907 ^ n31456 ;
  assign n31909 = n31908 ^ n31885 ;
  assign n31910 = n31906 & n31909 ;
  assign n31911 = n31910 ^ n31907 ;
  assign n31883 = n31352 ^ n31338 ;
  assign n32035 = n31911 ^ n31883 ;
  assign n32036 = ~n30601 & n32035 ;
  assign n32037 = n32036 ^ n31456 ;
  assign n31934 = n31903 ^ n31886 ;
  assign n31935 = ~n30580 & n31934 ;
  assign n31936 = n31935 ^ n31413 ;
  assign n31937 = n31936 ^ n30013 ;
  assign n31943 = n30404 & ~n31942 ;
  assign n31944 = n31943 ^ n31024 ;
  assign n31945 = n31944 ^ n30000 ;
  assign n32014 = ~n30428 & ~n31859 ;
  assign n32015 = n32014 ^ n31354 ;
  assign n31946 = n30435 & n31864 ;
  assign n31947 = n31946 ^ n31324 ;
  assign n31948 = n31947 ^ n29884 ;
  assign n31997 = ~n30438 & ~n31866 ;
  assign n31998 = n31997 ^ n31312 ;
  assign n31949 = n31843 ^ n31813 ;
  assign n31950 = ~n30552 & ~n31949 ;
  assign n31951 = n31950 ^ n31293 ;
  assign n31952 = n31951 ^ n29891 ;
  assign n31986 = n31840 ^ n31815 ;
  assign n31987 = n30440 & n31986 ;
  assign n31988 = n31987 ^ n31282 ;
  assign n31953 = n30540 & ~n31872 ;
  assign n31954 = n31953 ^ n31262 ;
  assign n31955 = n31954 ^ n29967 ;
  assign n31958 = ~n30533 & n31957 ;
  assign n31959 = n31958 ^ n31246 ;
  assign n31960 = n31959 ^ n30269 ;
  assign n31977 = n31976 ^ n31962 ;
  assign n31978 = ~n31963 & n31977 ;
  assign n31979 = n31978 ^ n29900 ;
  assign n31980 = n31979 ^ n31959 ;
  assign n31981 = n31960 & n31980 ;
  assign n31982 = n31981 ^ n30269 ;
  assign n31983 = n31982 ^ n31954 ;
  assign n31984 = n31955 & ~n31983 ;
  assign n31985 = n31984 ^ n29967 ;
  assign n31989 = n31988 ^ n31985 ;
  assign n31990 = n31951 ^ n29811 ;
  assign n31991 = n31990 ^ n31951 ;
  assign n31992 = n31991 ^ n31985 ;
  assign n31993 = n31989 & ~n31992 ;
  assign n31994 = n31993 ^ n31990 ;
  assign n31995 = n31952 & ~n31994 ;
  assign n31996 = n31995 ^ n29891 ;
  assign n31999 = n31998 ^ n31996 ;
  assign n32000 = n31947 ^ n29806 ;
  assign n32001 = n32000 ^ n31947 ;
  assign n32002 = n32001 ^ n31996 ;
  assign n32003 = ~n31999 & ~n32002 ;
  assign n32004 = n32003 ^ n32000 ;
  assign n32005 = n31948 & n32004 ;
  assign n32006 = n32005 ^ n29884 ;
  assign n32007 = n32006 ^ n30388 ;
  assign n32008 = n31855 ^ n31807 ;
  assign n32009 = n30432 & n32008 ;
  assign n32010 = n32009 ^ n31339 ;
  assign n32011 = n32010 ^ n32006 ;
  assign n32012 = n32007 & n32011 ;
  assign n32013 = n32012 ^ n30388 ;
  assign n32016 = n32015 ^ n32013 ;
  assign n32017 = n31944 ^ n30390 ;
  assign n32018 = n32017 ^ n32013 ;
  assign n32019 = n32018 ^ n31944 ;
  assign n32020 = n32016 & ~n32019 ;
  assign n32021 = n32020 ^ n32017 ;
  assign n32022 = n31945 & ~n32021 ;
  assign n32023 = n32022 ^ n30000 ;
  assign n31940 = n30573 & n31939 ;
  assign n31941 = n31940 ^ n31390 ;
  assign n32024 = n32023 ^ n31941 ;
  assign n32025 = n32023 ^ n30004 ;
  assign n32026 = ~n32024 & n32025 ;
  assign n32027 = n32026 ^ n30004 ;
  assign n32028 = n32027 ^ n31936 ;
  assign n32029 = n31937 & ~n32028 ;
  assign n32030 = n32029 ^ n30013 ;
  assign n31930 = n31885 ^ n31442 ;
  assign n31931 = n31930 ^ n31905 ;
  assign n31932 = n30424 & n31931 ;
  assign n31933 = n31932 ^ n31442 ;
  assign n32031 = n32030 ^ n31933 ;
  assign n32032 = n32030 ^ n30408 ;
  assign n32033 = n32031 & ~n32032 ;
  assign n32034 = n32033 ^ n30408 ;
  assign n32038 = n32037 ^ n32034 ;
  assign n32039 = n32037 ^ n30030 ;
  assign n32040 = ~n32038 & n32039 ;
  assign n32041 = n32040 ^ n30030 ;
  assign n31882 = n31367 ^ n31353 ;
  assign n31925 = n31882 ^ n31483 ;
  assign n31884 = n31883 ^ n31456 ;
  assign n31912 = ~n31884 & n31911 ;
  assign n31913 = n31912 ^ n31456 ;
  assign n31926 = n31925 ^ n31913 ;
  assign n31927 = ~n30611 & n31926 ;
  assign n31928 = n31927 ^ n31483 ;
  assign n31929 = n31928 ^ n29876 ;
  assign n32164 = n32041 ^ n31929 ;
  assign n32076 = n31933 ^ n30408 ;
  assign n32077 = n32076 ^ n32030 ;
  assign n32078 = n32077 ^ x253 ;
  assign n32149 = n32027 ^ n31937 ;
  assign n32079 = n32021 ^ n30000 ;
  assign n32080 = n32079 ^ x240 ;
  assign n32083 = n32010 ^ n32007 ;
  assign n32084 = n32083 ^ x242 ;
  assign n32085 = n32004 ^ n29884 ;
  assign n32086 = n32085 ^ x243 ;
  assign n32087 = n31996 ^ n29806 ;
  assign n32088 = n32087 ^ n31998 ;
  assign n32089 = n32088 ^ x244 ;
  assign n32090 = n31994 ^ n29891 ;
  assign n32091 = n32090 ^ x245 ;
  assign n32117 = n31988 ^ n29811 ;
  assign n32118 = n32117 ^ n31985 ;
  assign n32092 = n31982 ^ n29967 ;
  assign n32093 = n32092 ^ n31954 ;
  assign n32094 = n32093 ^ x247 ;
  assign n32108 = n31979 ^ n31960 ;
  assign n32096 = n32095 ^ x233 ;
  assign n32105 = n32104 ^ n32095 ;
  assign n32106 = n32096 & ~n32105 ;
  assign n32107 = n32106 ^ x233 ;
  assign n32109 = n32108 ^ n32107 ;
  assign n32110 = n32093 ^ x232 ;
  assign n32111 = n32110 ^ n32093 ;
  assign n32112 = n32111 ^ n32107 ;
  assign n32113 = n32109 & n32112 ;
  assign n32114 = n32113 ^ n32110 ;
  assign n32115 = n32094 & ~n32114 ;
  assign n32116 = n32115 ^ x247 ;
  assign n32119 = n32118 ^ n32116 ;
  assign n32120 = n32090 ^ x246 ;
  assign n32121 = n32120 ^ n32090 ;
  assign n32122 = n32121 ^ n32116 ;
  assign n32123 = ~n32119 & n32122 ;
  assign n32124 = n32123 ^ n32120 ;
  assign n32125 = ~n32091 & n32124 ;
  assign n32126 = n32125 ^ x245 ;
  assign n32127 = n32126 ^ n32088 ;
  assign n32128 = n32089 & ~n32127 ;
  assign n32129 = n32128 ^ x244 ;
  assign n32130 = n32129 ^ n32085 ;
  assign n32131 = n32086 & ~n32130 ;
  assign n32132 = n32131 ^ x243 ;
  assign n32133 = n32132 ^ n32083 ;
  assign n32134 = n32084 & ~n32133 ;
  assign n32135 = n32134 ^ x242 ;
  assign n32081 = n32015 ^ n30390 ;
  assign n32082 = n32081 ^ n32013 ;
  assign n32136 = n32135 ^ n32082 ;
  assign n32137 = n32135 ^ x241 ;
  assign n32138 = n32136 & n32137 ;
  assign n32139 = n32138 ^ x241 ;
  assign n32140 = n32139 ^ n32079 ;
  assign n32141 = n32080 & ~n32140 ;
  assign n32142 = n32141 ^ x240 ;
  assign n32143 = n32142 ^ x255 ;
  assign n32144 = n31941 ^ n30004 ;
  assign n32145 = n32144 ^ n32023 ;
  assign n32146 = n32145 ^ n32142 ;
  assign n32147 = n32143 & ~n32146 ;
  assign n32148 = n32147 ^ x255 ;
  assign n32150 = n32149 ^ n32148 ;
  assign n32151 = n32077 ^ x254 ;
  assign n32152 = n32151 ^ n32148 ;
  assign n32153 = n32152 ^ n32077 ;
  assign n32154 = ~n32150 & n32153 ;
  assign n32155 = n32154 ^ n32151 ;
  assign n32156 = n32078 & ~n32155 ;
  assign n32157 = n32156 ^ x253 ;
  assign n32158 = n32157 ^ x252 ;
  assign n32159 = n32034 ^ n30030 ;
  assign n32160 = n32159 ^ n32037 ;
  assign n32161 = n32160 ^ n32157 ;
  assign n32162 = n32158 & n32161 ;
  assign n32163 = n32162 ^ x252 ;
  assign n32165 = n32164 ^ n32163 ;
  assign n32042 = n32041 ^ n31928 ;
  assign n32043 = n31929 & n32042 ;
  assign n32044 = n32043 ^ n29876 ;
  assign n32166 = n32044 ^ n30621 ;
  assign n31920 = n31382 ^ n31368 ;
  assign n31914 = n31913 ^ n31882 ;
  assign n31915 = n31503 ^ n31483 ;
  assign n31916 = n31915 ^ n31503 ;
  assign n31917 = n31916 ^ n31882 ;
  assign n31918 = ~n31914 & ~n31917 ;
  assign n31919 = n31918 ^ n31915 ;
  assign n31921 = n31920 ^ n31919 ;
  assign n31922 = ~n30624 & ~n31921 ;
  assign n31923 = n31922 ^ n31503 ;
  assign n32167 = n32166 ^ n31923 ;
  assign n32168 = n32167 ^ x251 ;
  assign n32169 = n32168 ^ n32163 ;
  assign n32170 = n32169 ^ n32167 ;
  assign n32171 = n32165 & n32170 ;
  assign n32172 = n32171 ^ n32168 ;
  assign n32181 = n32172 ^ x250 ;
  assign n32182 = n32164 ^ x251 ;
  assign n32183 = n32182 ^ n32163 ;
  assign n32184 = n32160 ^ n32158 ;
  assign n32185 = n32155 ^ x253 ;
  assign n32186 = n32149 ^ x254 ;
  assign n32187 = n32186 ^ n32148 ;
  assign n32188 = n32145 ^ n32143 ;
  assign n32189 = n32139 ^ n32080 ;
  assign n32190 = n32082 ^ x241 ;
  assign n32191 = n32190 ^ n32135 ;
  assign n32198 = n32195 & ~n32197 ;
  assign n32199 = n32107 ^ x232 ;
  assign n32200 = n32199 ^ n32108 ;
  assign n32201 = n32198 & n32200 ;
  assign n32202 = n32114 ^ x247 ;
  assign n32203 = ~n32201 & n32202 ;
  assign n32204 = n32118 ^ x246 ;
  assign n32205 = n32204 ^ n32116 ;
  assign n32206 = ~n32203 & ~n32205 ;
  assign n32207 = n32124 ^ x245 ;
  assign n32208 = ~n32206 & ~n32207 ;
  assign n32209 = n32126 ^ n32089 ;
  assign n32210 = ~n32208 & ~n32209 ;
  assign n32211 = n32129 ^ n32086 ;
  assign n32212 = ~n32210 & n32211 ;
  assign n32213 = n32132 ^ x242 ;
  assign n32214 = n32213 ^ n32083 ;
  assign n32215 = ~n32212 & ~n32214 ;
  assign n32216 = ~n32191 & ~n32215 ;
  assign n32217 = n32189 & n32216 ;
  assign n32218 = ~n32188 & ~n32217 ;
  assign n32219 = ~n32187 & n32218 ;
  assign n32220 = n32185 & ~n32219 ;
  assign n32221 = ~n32184 & n32220 ;
  assign n32222 = ~n32183 & n32221 ;
  assign n32223 = n32181 & n32222 ;
  assign n31924 = n31923 ^ n30621 ;
  assign n32045 = n32044 ^ n31923 ;
  assign n32046 = n31924 & n32045 ;
  assign n32047 = n32046 ^ n30621 ;
  assign n32073 = n32047 ^ n30633 ;
  assign n32048 = n31404 ^ n31383 ;
  assign n32050 = n32048 ^ n31503 ;
  assign n32049 = n32048 ^ n31920 ;
  assign n32051 = n32050 ^ n32049 ;
  assign n32052 = ~n31919 & ~n32051 ;
  assign n32053 = n32052 ^ n32050 ;
  assign n32054 = n32053 ^ n31525 ;
  assign n32055 = n30636 & n32054 ;
  assign n32056 = n32055 ^ n31525 ;
  assign n32074 = n32073 ^ n32056 ;
  assign n32174 = n32074 ^ x250 ;
  assign n32173 = n32167 ^ n32074 ;
  assign n32175 = n32174 ^ n32173 ;
  assign n32176 = ~n32172 & n32175 ;
  assign n32177 = n32176 ^ n32174 ;
  assign n32180 = n32177 ^ x249 ;
  assign n32226 = n32223 ^ n32180 ;
  assign n32227 = n32226 ^ n31602 ;
  assign n32257 = n32221 ^ n32183 ;
  assign n32228 = n32220 ^ n32184 ;
  assign n32229 = n32228 ^ n31610 ;
  assign n32231 = n32218 ^ n32187 ;
  assign n32232 = n32231 ^ n31618 ;
  assign n32240 = n32217 ^ n32188 ;
  assign n32235 = n32216 ^ n32189 ;
  assign n32233 = n32215 ^ n32191 ;
  assign n32234 = n31628 & n32233 ;
  assign n32236 = n32235 ^ n32234 ;
  assign n32237 = n32235 ^ n31625 ;
  assign n32238 = ~n32236 & n32237 ;
  assign n32239 = n32238 ^ n31625 ;
  assign n32241 = n32240 ^ n32239 ;
  assign n32242 = n32231 ^ n31622 ;
  assign n32243 = n32242 ^ n32231 ;
  assign n32244 = n32243 ^ n32239 ;
  assign n32245 = n32241 & ~n32244 ;
  assign n32246 = n32245 ^ n32242 ;
  assign n32247 = n32232 & n32246 ;
  assign n32248 = n32247 ^ n31618 ;
  assign n32230 = n32219 ^ n32185 ;
  assign n32249 = n32248 ^ n32230 ;
  assign n32250 = n32228 ^ n31614 ;
  assign n32251 = n32250 ^ n32230 ;
  assign n32252 = n32251 ^ n32228 ;
  assign n32253 = n32249 & ~n32252 ;
  assign n32254 = n32253 ^ n32250 ;
  assign n32255 = ~n32229 & n32254 ;
  assign n32256 = n32255 ^ n31610 ;
  assign n32258 = n32257 ^ n32256 ;
  assign n32259 = n32222 ^ n32181 ;
  assign n32260 = n32259 ^ n31606 ;
  assign n32261 = n32260 ^ n32256 ;
  assign n32262 = n32261 ^ n32259 ;
  assign n32263 = n32258 & n32262 ;
  assign n32264 = n32263 ^ n32260 ;
  assign n32266 = n32226 ^ n31654 ;
  assign n32265 = n32259 ^ n32226 ;
  assign n32267 = n32266 ^ n32265 ;
  assign n32268 = ~n32264 & n32267 ;
  assign n32269 = n32268 ^ n32266 ;
  assign n32270 = n32227 & ~n32269 ;
  assign n32271 = n32270 ^ n31602 ;
  assign n32224 = n32180 & ~n32223 ;
  assign n32075 = n32074 ^ x249 ;
  assign n32178 = ~n32075 & n32177 ;
  assign n32067 = n32048 ^ n31525 ;
  assign n32068 = n32053 & ~n32067 ;
  assign n32064 = n31426 ^ n31405 ;
  assign n32065 = n32064 ^ n31571 ;
  assign n32066 = n32065 ^ n32048 ;
  assign n32069 = n32068 ^ n32066 ;
  assign n32070 = ~n30646 & n32069 ;
  assign n32062 = x249 ^ x248 ;
  assign n32060 = n30633 ^ n30196 ;
  assign n32061 = n32060 ^ n31571 ;
  assign n32063 = n32062 ^ n32061 ;
  assign n32071 = n32070 ^ n32063 ;
  assign n32057 = n32056 ^ n32047 ;
  assign n32058 = n32056 ^ n30633 ;
  assign n32059 = n32057 & n32058 ;
  assign n32072 = n32071 ^ n32059 ;
  assign n32179 = n32178 ^ n32072 ;
  assign n32225 = n32224 ^ n32179 ;
  assign n32272 = n32271 ^ n32225 ;
  assign n32273 = n32271 ^ n31599 ;
  assign n32274 = n32272 & ~n32273 ;
  assign n32275 = n32274 ^ n31599 ;
  assign n32276 = n32275 ^ n31777 ;
  assign n32277 = ~n31881 & n32276 ;
  assign n32278 = n32277 ^ n31672 ;
  assign n32280 = n32279 ^ n32278 ;
  assign n32281 = n31879 ^ n31745 ;
  assign n32282 = n32281 ^ n31879 ;
  assign n32283 = n32282 ^ n32278 ;
  assign n32284 = ~n32280 & ~n32283 ;
  assign n32285 = n32284 ^ n32281 ;
  assign n32286 = ~n31880 & n32285 ;
  assign n32287 = n32286 ^ n31766 ;
  assign n31878 = n31785 ^ n31783 ;
  assign n32288 = n32287 ^ n31878 ;
  assign n32289 = n32287 ^ n31965 ;
  assign n32290 = n32288 & n32289 ;
  assign n32291 = n32290 ^ n31965 ;
  assign n32292 = n32291 ^ n31875 ;
  assign n32293 = ~n31877 & ~n32292 ;
  assign n32294 = n32293 ^ n31876 ;
  assign n31874 = n31788 ^ n31787 ;
  assign n32295 = n32294 ^ n31874 ;
  assign n32296 = n32294 ^ n31957 ;
  assign n32297 = n32295 & n32296 ;
  assign n32299 = n32298 ^ n32297 ;
  assign n32300 = ~n31873 & ~n32299 ;
  assign n32301 = n32300 ^ n31872 ;
  assign n31870 = n31793 ^ n31792 ;
  assign n32302 = n32301 ^ n31870 ;
  assign n32303 = n31796 ^ n31794 ;
  assign n32304 = n32303 ^ n31986 ;
  assign n32305 = n32304 ^ n31870 ;
  assign n32306 = n32305 ^ n32303 ;
  assign n32307 = n32302 & n32306 ;
  assign n32308 = n32307 ^ n32304 ;
  assign n32310 = n31949 ^ n31868 ;
  assign n32309 = n32303 ^ n31868 ;
  assign n32311 = n32310 ^ n32309 ;
  assign n32312 = n32308 & n32311 ;
  assign n32313 = n32312 ^ n32310 ;
  assign n32314 = n31869 & ~n32313 ;
  assign n31867 = n31866 ^ n31864 ;
  assign n32315 = n32314 ^ n31867 ;
  assign n32316 = ~n31865 & ~n32315 ;
  assign n32317 = n32316 ^ n31864 ;
  assign n31861 = n31803 ^ n31802 ;
  assign n32318 = n32317 ^ n31861 ;
  assign n32319 = n32317 ^ n32008 ;
  assign n32320 = ~n32318 & n32319 ;
  assign n32321 = n32320 ^ n32008 ;
  assign n32322 = n32321 ^ n31805 ;
  assign n32323 = ~n31860 & ~n32322 ;
  assign n32324 = n32323 ^ n31859 ;
  assign n32703 = n32325 ^ n32324 ;
  assign n32704 = n32326 & ~n32703 ;
  assign n32705 = n32704 ^ n31942 ;
  assign n32708 = n32707 ^ n32705 ;
  assign n32345 = n31957 ^ n31874 ;
  assign n32346 = n32345 ^ n32294 ;
  assign n32347 = ~n31246 & ~n32346 ;
  assign n32348 = n32347 ^ n31957 ;
  assign n32517 = n32348 ^ n30533 ;
  assign n32349 = n32291 ^ n31877 ;
  assign n32350 = ~n31232 & n32349 ;
  assign n32351 = n32350 ^ n31876 ;
  assign n32352 = n32351 ^ n30444 ;
  assign n32449 = n31965 ^ n31878 ;
  assign n32450 = n32449 ^ n32287 ;
  assign n32451 = n31217 & n32450 ;
  assign n32452 = n32451 ^ n31965 ;
  assign n32353 = n32285 ^ n31766 ;
  assign n32354 = n31200 & n32353 ;
  assign n32355 = n32354 ^ n31766 ;
  assign n32356 = n32355 ^ n30450 ;
  assign n32361 = n32225 ^ n31599 ;
  assign n32362 = n32361 ^ n32271 ;
  assign n32363 = n31151 & ~n32362 ;
  assign n32364 = n32363 ^ n31599 ;
  assign n32365 = n32364 ^ n30510 ;
  assign n32369 = n32264 ^ n31654 ;
  assign n32370 = ~n31118 & ~n32369 ;
  assign n32371 = n32370 ^ n31654 ;
  assign n32372 = n32371 ^ n30460 ;
  assign n32377 = n32254 ^ n31610 ;
  assign n32378 = n31088 & n32377 ;
  assign n32379 = n32378 ^ n31610 ;
  assign n32380 = n32379 ^ n30465 ;
  assign n32385 = n32246 ^ n31618 ;
  assign n32386 = ~n31060 & n32385 ;
  assign n32387 = n32386 ^ n31618 ;
  assign n32388 = n32387 ^ n30471 ;
  assign n32402 = n32239 ^ n31622 ;
  assign n32403 = n32402 ^ n32240 ;
  assign n32404 = ~n31049 & ~n32403 ;
  assign n32405 = n32404 ^ n31622 ;
  assign n32394 = n32234 ^ n31625 ;
  assign n32395 = n32394 ^ n32235 ;
  assign n32396 = ~n31034 & ~n32395 ;
  assign n32397 = n32396 ^ n31625 ;
  assign n32389 = n32233 ^ n31538 ;
  assign n32390 = n32389 ^ n31026 ;
  assign n32391 = ~n31026 & ~n32390 ;
  assign n32392 = n32391 ^ n31628 ;
  assign n32393 = n30925 & ~n32392 ;
  assign n32398 = n32397 ^ n32393 ;
  assign n32399 = n32397 ^ n30479 ;
  assign n32400 = n32398 & ~n32399 ;
  assign n32401 = n32400 ^ n30479 ;
  assign n32406 = n32405 ^ n32401 ;
  assign n32407 = n32387 ^ n30474 ;
  assign n32408 = n32407 ^ n32387 ;
  assign n32409 = n32408 ^ n32401 ;
  assign n32410 = ~n32406 & ~n32409 ;
  assign n32411 = n32410 ^ n32407 ;
  assign n32412 = n32388 & ~n32411 ;
  assign n32413 = n32412 ^ n30471 ;
  assign n32381 = n32248 ^ n31614 ;
  assign n32382 = n32381 ^ n32230 ;
  assign n32383 = ~n31071 & n32382 ;
  assign n32384 = n32383 ^ n31614 ;
  assign n32414 = n32413 ^ n32384 ;
  assign n32415 = n32413 ^ n30468 ;
  assign n32416 = ~n32414 & n32415 ;
  assign n32417 = n32416 ^ n30468 ;
  assign n32418 = n32417 ^ n32379 ;
  assign n32419 = n32380 & ~n32418 ;
  assign n32420 = n32419 ^ n30465 ;
  assign n32373 = n32257 ^ n31606 ;
  assign n32374 = n32373 ^ n32256 ;
  assign n32375 = ~n31030 & n32374 ;
  assign n32376 = n32375 ^ n31606 ;
  assign n32421 = n32420 ^ n32376 ;
  assign n32422 = n32420 ^ n30462 ;
  assign n32423 = ~n32421 & n32422 ;
  assign n32424 = n32423 ^ n30462 ;
  assign n32425 = n32424 ^ n32371 ;
  assign n32426 = ~n32372 & ~n32425 ;
  assign n32427 = n32426 ^ n30460 ;
  assign n32366 = n32269 ^ n31602 ;
  assign n32367 = n31136 & ~n32366 ;
  assign n32368 = n32367 ^ n31602 ;
  assign n32428 = n32427 ^ n32368 ;
  assign n32429 = n32427 ^ n30457 ;
  assign n32430 = n32428 & n32429 ;
  assign n32431 = n32430 ^ n30457 ;
  assign n32432 = n32431 ^ n32364 ;
  assign n32433 = ~n32365 & ~n32432 ;
  assign n32434 = n32433 ^ n30510 ;
  assign n32435 = n32434 ^ n30455 ;
  assign n32438 = n32434 ^ n31671 ;
  assign n32436 = n32275 ^ n31881 ;
  assign n32437 = n31165 & n32436 ;
  assign n32439 = n32438 ^ n32437 ;
  assign n32440 = n32435 & n32439 ;
  assign n32441 = n32440 ^ n30455 ;
  assign n32357 = n32279 ^ n31745 ;
  assign n32358 = n32357 ^ n32278 ;
  assign n32359 = ~n31185 & ~n32358 ;
  assign n32360 = n32359 ^ n31745 ;
  assign n32442 = n32441 ^ n32360 ;
  assign n32443 = n32441 ^ n30452 ;
  assign n32444 = ~n32442 & n32443 ;
  assign n32445 = n32444 ^ n30452 ;
  assign n32446 = n32445 ^ n32355 ;
  assign n32447 = ~n32356 & ~n32446 ;
  assign n32448 = n32447 ^ n30450 ;
  assign n32453 = n32452 ^ n32448 ;
  assign n32454 = n32351 ^ n30446 ;
  assign n32455 = n32454 ^ n32448 ;
  assign n32456 = n32455 ^ n32351 ;
  assign n32457 = n32453 & n32456 ;
  assign n32458 = n32457 ^ n32454 ;
  assign n32459 = n32352 & ~n32458 ;
  assign n32460 = n32459 ^ n30444 ;
  assign n32518 = n32517 ^ n32460 ;
  assign n32519 = n32518 ^ x456 ;
  assign n32601 = n32458 ^ n30444 ;
  assign n32520 = n32452 ^ n30446 ;
  assign n32521 = n32520 ^ n32448 ;
  assign n32522 = n32521 ^ x458 ;
  assign n32525 = n32360 ^ n30452 ;
  assign n32526 = n32525 ^ n32441 ;
  assign n32527 = n32526 ^ x460 ;
  assign n32529 = n32431 ^ n32365 ;
  assign n32530 = n32529 ^ x462 ;
  assign n32570 = n32424 ^ n32372 ;
  assign n32533 = n32417 ^ n30465 ;
  assign n32534 = n32533 ^ n32379 ;
  assign n32535 = n32534 ^ x450 ;
  assign n32536 = n32384 ^ n30468 ;
  assign n32537 = n32536 ^ n32413 ;
  assign n32538 = n32537 ^ x451 ;
  assign n32554 = n32411 ^ n30471 ;
  assign n32548 = n32405 ^ n30474 ;
  assign n32549 = n32548 ^ n32401 ;
  assign n32542 = n32393 ^ n30479 ;
  assign n32543 = n32542 ^ n32397 ;
  assign n32539 = n31538 ^ n30926 ;
  assign n32540 = n32539 ^ n32391 ;
  assign n32541 = x455 & ~n32540 ;
  assign n32544 = n32543 ^ n32541 ;
  assign n32545 = n32543 ^ x454 ;
  assign n32546 = n32544 & ~n32545 ;
  assign n32547 = n32546 ^ x454 ;
  assign n32550 = n32549 ^ n32547 ;
  assign n32551 = n32549 ^ x453 ;
  assign n32552 = n32550 & ~n32551 ;
  assign n32553 = n32552 ^ x453 ;
  assign n32555 = n32554 ^ n32553 ;
  assign n32556 = n32537 ^ x452 ;
  assign n32557 = n32556 ^ n32537 ;
  assign n32558 = n32557 ^ n32553 ;
  assign n32559 = n32555 & n32558 ;
  assign n32560 = n32559 ^ n32556 ;
  assign n32561 = ~n32538 & n32560 ;
  assign n32562 = n32561 ^ x451 ;
  assign n32563 = n32562 ^ n32534 ;
  assign n32564 = ~n32535 & n32563 ;
  assign n32565 = n32564 ^ x450 ;
  assign n32531 = n32376 ^ n30462 ;
  assign n32532 = n32531 ^ n32420 ;
  assign n32566 = n32565 ^ n32532 ;
  assign n32567 = n32565 ^ x449 ;
  assign n32568 = n32566 & n32567 ;
  assign n32569 = n32568 ^ x449 ;
  assign n32571 = n32570 ^ n32569 ;
  assign n32572 = n32368 ^ n30457 ;
  assign n32573 = n32572 ^ n32427 ;
  assign n32574 = n32573 ^ x448 ;
  assign n32575 = n32574 ^ n32573 ;
  assign n32576 = n32575 ^ n32569 ;
  assign n32577 = ~n32571 & n32576 ;
  assign n32578 = n32577 ^ n32574 ;
  assign n32580 = n32529 ^ x463 ;
  assign n32579 = n32573 ^ n32529 ;
  assign n32581 = n32580 ^ n32579 ;
  assign n32582 = n32578 & ~n32581 ;
  assign n32583 = n32582 ^ n32580 ;
  assign n32584 = ~n32530 & n32583 ;
  assign n32585 = n32584 ^ x462 ;
  assign n32528 = n32439 ^ n30455 ;
  assign n32586 = n32585 ^ n32528 ;
  assign n32587 = n32585 ^ x461 ;
  assign n32588 = ~n32586 & n32587 ;
  assign n32589 = n32588 ^ x461 ;
  assign n32590 = n32589 ^ n32526 ;
  assign n32591 = ~n32527 & n32590 ;
  assign n32592 = n32591 ^ x460 ;
  assign n32523 = n32445 ^ n30450 ;
  assign n32524 = n32523 ^ n32355 ;
  assign n32593 = n32592 ^ n32524 ;
  assign n32594 = n32521 ^ x459 ;
  assign n32595 = n32594 ^ n32524 ;
  assign n32596 = n32595 ^ n32521 ;
  assign n32597 = ~n32593 & n32596 ;
  assign n32598 = n32597 ^ n32594 ;
  assign n32599 = ~n32522 & n32598 ;
  assign n32600 = n32599 ^ x458 ;
  assign n32602 = n32601 ^ n32600 ;
  assign n32603 = n32518 ^ x457 ;
  assign n32604 = n32603 ^ n32600 ;
  assign n32605 = n32604 ^ n32518 ;
  assign n32606 = ~n32602 & n32605 ;
  assign n32607 = n32606 ^ n32603 ;
  assign n32608 = ~n32519 & n32607 ;
  assign n32609 = n32608 ^ x456 ;
  assign n32461 = n32460 ^ n32348 ;
  assign n32462 = n32460 ^ n30533 ;
  assign n32463 = ~n32461 & ~n32462 ;
  assign n32464 = n32463 ^ n30533 ;
  assign n32515 = n32464 ^ n30540 ;
  assign n32465 = n32299 ^ n31871 ;
  assign n32466 = ~n31262 & ~n32465 ;
  assign n32467 = n32466 ^ n31872 ;
  assign n32516 = n32515 ^ n32467 ;
  assign n32610 = n32609 ^ n32516 ;
  assign n32611 = n32609 ^ x471 ;
  assign n32612 = ~n32610 & n32611 ;
  assign n32613 = n32612 ^ x471 ;
  assign n32684 = n32613 ^ x470 ;
  assign n32468 = n32467 ^ n32464 ;
  assign n32469 = n32467 ^ n30540 ;
  assign n32470 = ~n32468 & ~n32469 ;
  assign n32471 = n32470 ^ n30540 ;
  assign n32340 = n31986 ^ n31870 ;
  assign n32341 = n32340 ^ n32301 ;
  assign n32342 = n31282 & ~n32341 ;
  assign n32343 = n32342 ^ n31986 ;
  assign n32344 = n32343 ^ n30440 ;
  assign n32614 = n32471 ^ n32344 ;
  assign n32685 = n32684 ^ n32614 ;
  assign n32641 = n32540 ^ x455 ;
  assign n32642 = n32541 ^ x454 ;
  assign n32643 = n32642 ^ n32543 ;
  assign n32644 = n32641 & n32643 ;
  assign n32645 = n32547 ^ x453 ;
  assign n32646 = n32645 ^ n32549 ;
  assign n32647 = n32644 & n32646 ;
  assign n32648 = n32554 ^ x452 ;
  assign n32649 = n32648 ^ n32553 ;
  assign n32650 = ~n32647 & ~n32649 ;
  assign n32651 = n32560 ^ x451 ;
  assign n32652 = n32650 & ~n32651 ;
  assign n32653 = n32562 ^ n32535 ;
  assign n32654 = ~n32652 & n32653 ;
  assign n32655 = n32532 ^ x449 ;
  assign n32656 = n32655 ^ n32565 ;
  assign n32657 = ~n32654 & ~n32656 ;
  assign n32658 = n32570 ^ x448 ;
  assign n32659 = n32658 ^ n32569 ;
  assign n32660 = ~n32657 & ~n32659 ;
  assign n32661 = n32578 ^ x463 ;
  assign n32662 = n32660 & n32661 ;
  assign n32663 = n32583 ^ x462 ;
  assign n32664 = n32662 & n32663 ;
  assign n32665 = n32528 ^ x461 ;
  assign n32666 = n32665 ^ n32585 ;
  assign n32667 = ~n32664 & n32666 ;
  assign n32668 = n32589 ^ x460 ;
  assign n32669 = n32668 ^ n32526 ;
  assign n32670 = n32667 & ~n32669 ;
  assign n32671 = n32592 ^ x459 ;
  assign n32672 = n32671 ^ n32524 ;
  assign n32673 = n32670 & n32672 ;
  assign n32674 = n32598 ^ x458 ;
  assign n32675 = ~n32673 & n32674 ;
  assign n32676 = n32601 ^ x457 ;
  assign n32677 = n32676 ^ n32600 ;
  assign n32678 = ~n32675 & n32677 ;
  assign n32679 = n32607 ^ x456 ;
  assign n32680 = n32678 & ~n32679 ;
  assign n32681 = n32516 ^ x471 ;
  assign n32682 = n32681 ^ n32609 ;
  assign n32683 = n32680 & n32682 ;
  assign n32719 = n32685 ^ n32683 ;
  assign n32802 = n32719 ^ n32390 ;
  assign n32811 = n31628 & ~n32802 ;
  assign n32812 = n32811 ^ n32389 ;
  assign n32997 = n32812 ^ x167 ;
  assign n32916 = x167 & n32812 ;
  assign n32918 = n32916 ^ x166 ;
  assign n32615 = n32614 ^ n32613 ;
  assign n32616 = n32614 ^ x470 ;
  assign n32617 = ~n32615 & n32616 ;
  assign n32618 = n32617 ^ x470 ;
  assign n32472 = n32471 ^ n32343 ;
  assign n32473 = n32344 & ~n32472 ;
  assign n32474 = n32473 ^ n30440 ;
  assign n32512 = n32474 ^ n30552 ;
  assign n32475 = n32308 ^ n31949 ;
  assign n32476 = n31293 & n32475 ;
  assign n32477 = n32476 ^ n31949 ;
  assign n32513 = n32512 ^ n32477 ;
  assign n32514 = n32513 ^ x469 ;
  assign n32687 = n32618 ^ n32514 ;
  assign n32686 = n32683 & n32685 ;
  assign n32722 = n32687 ^ n32686 ;
  assign n32720 = n32390 & n32719 ;
  assign n32721 = n32720 ^ n32395 ;
  assign n32815 = n32722 ^ n32721 ;
  assign n32816 = n31625 & n32815 ;
  assign n32817 = n32816 ^ n32395 ;
  assign n32813 = ~n31026 & ~n32812 ;
  assign n32814 = n32813 ^ n31034 ;
  assign n32915 = n32817 ^ n32814 ;
  assign n32998 = n32918 ^ n32915 ;
  assign n32999 = n32997 & n32998 ;
  assign n32478 = n32477 ^ n32474 ;
  assign n32336 = n32313 ^ n31866 ;
  assign n32337 = n31312 & ~n32336 ;
  assign n32338 = n32337 ^ n31866 ;
  assign n32479 = n32338 ^ n30552 ;
  assign n32480 = n32479 ^ n32474 ;
  assign n32481 = n32480 ^ n32338 ;
  assign n32482 = n32478 & ~n32481 ;
  assign n32483 = n32482 ^ n32479 ;
  assign n32511 = n32483 ^ n30438 ;
  assign n32689 = n32511 ^ x468 ;
  assign n32619 = n32618 ^ n32513 ;
  assign n32620 = n32514 & ~n32619 ;
  assign n32621 = n32620 ^ x469 ;
  assign n32690 = n32689 ^ n32621 ;
  assign n32688 = ~n32686 & ~n32687 ;
  assign n32718 = n32690 ^ n32688 ;
  assign n32807 = n32718 ^ n32403 ;
  assign n32723 = n32722 ^ n32720 ;
  assign n32724 = n32721 & n32723 ;
  assign n32725 = n32724 ^ n32395 ;
  assign n32808 = n32807 ^ n32725 ;
  assign n32809 = ~n31622 & ~n32808 ;
  assign n32810 = n32809 ^ n32403 ;
  assign n32913 = n32810 ^ n31049 ;
  assign n32818 = n32817 ^ n32813 ;
  assign n32819 = ~n32814 & n32818 ;
  assign n32820 = n32819 ^ n31034 ;
  assign n32914 = n32913 ^ n32820 ;
  assign n32995 = n32914 ^ x165 ;
  assign n32917 = n32916 ^ n32915 ;
  assign n32919 = ~n32917 & n32918 ;
  assign n32920 = n32919 ^ x166 ;
  assign n32996 = n32995 ^ n32920 ;
  assign n33400 = n32999 ^ n32996 ;
  assign n33369 = n32661 ^ n32660 ;
  assign n32498 = n32321 ^ n31860 ;
  assign n32327 = n32326 ^ n32324 ;
  assign n33367 = n32498 ^ n32327 ;
  assign n33363 = n32659 ^ n32657 ;
  assign n33350 = n32656 ^ n32654 ;
  assign n32331 = n32008 ^ n31861 ;
  assign n32332 = n32331 ^ n32317 ;
  assign n33351 = n33350 ^ n32332 ;
  assign n33352 = n32653 ^ n32652 ;
  assign n32486 = n32315 ^ n31862 ;
  assign n33353 = n33352 ^ n32486 ;
  assign n33083 = n32211 ^ n32210 ;
  assign n32873 = n32205 ^ n32203 ;
  assign n32874 = n32873 ^ n32035 ;
  assign n32757 = n32706 ^ n32705 ;
  assign n32760 = n32705 ^ n31939 ;
  assign n32761 = ~n32757 & ~n32760 ;
  assign n32758 = n31939 ^ n31934 ;
  assign n32762 = n32761 ^ n32758 ;
  assign n32787 = n31934 ^ n31931 ;
  assign n32763 = n32200 ^ n32198 ;
  assign n32786 = n32763 ^ n31931 ;
  assign n32788 = n32787 ^ n32786 ;
  assign n32789 = n32762 & n32788 ;
  assign n32790 = n32789 ^ n32787 ;
  assign n32791 = n32202 ^ n32201 ;
  assign n32875 = n32791 ^ n31931 ;
  assign n32876 = n32790 & n32875 ;
  assign n32877 = n32876 ^ n31931 ;
  assign n32965 = n32877 ^ n32873 ;
  assign n32969 = n32874 & ~n32965 ;
  assign n32966 = n32035 ^ n31926 ;
  assign n32970 = n32969 ^ n32966 ;
  assign n32971 = n32207 ^ n32206 ;
  assign n33030 = n32971 ^ n31926 ;
  assign n33031 = n32970 & ~n33030 ;
  assign n33032 = n33031 ^ n31926 ;
  assign n33028 = n32209 ^ n32208 ;
  assign n33077 = n33032 ^ n33028 ;
  assign n33078 = n32054 ^ n31921 ;
  assign n33079 = n33078 ^ n32054 ;
  assign n33080 = n33079 ^ n33028 ;
  assign n33081 = ~n33077 & ~n33080 ;
  assign n33082 = n33081 ^ n33078 ;
  assign n33084 = n33083 ^ n33082 ;
  assign n33085 = ~n31525 & ~n33084 ;
  assign n33086 = n33085 ^ n32054 ;
  assign n33087 = n33086 ^ n30636 ;
  assign n33029 = n33028 ^ n31921 ;
  assign n33033 = n33032 ^ n33029 ;
  assign n33034 = n31503 & ~n33033 ;
  assign n33035 = n33034 ^ n31921 ;
  assign n32792 = n32791 ^ n32790 ;
  assign n32793 = n31442 & n32792 ;
  assign n32794 = n32793 ^ n31931 ;
  assign n32795 = n32794 ^ n30424 ;
  assign n32709 = ~n31390 & n32708 ;
  assign n32710 = n32709 ^ n31939 ;
  assign n32328 = ~n31024 & ~n32327 ;
  assign n32329 = n32328 ^ n31942 ;
  assign n32330 = n32329 ^ n30404 ;
  assign n32333 = ~n31339 & n32332 ;
  assign n32334 = n32333 ^ n32008 ;
  assign n32335 = n32334 ^ n30432 ;
  assign n32487 = n31324 & n32486 ;
  assign n32488 = n32487 ^ n31864 ;
  assign n32339 = n32338 ^ n30438 ;
  assign n32484 = n32339 & ~n32483 ;
  assign n32485 = n32484 ^ n30438 ;
  assign n32489 = n32488 ^ n32485 ;
  assign n32490 = n32334 ^ n30435 ;
  assign n32491 = n32490 ^ n32334 ;
  assign n32492 = n32491 ^ n32485 ;
  assign n32493 = n32489 & ~n32492 ;
  assign n32494 = n32493 ^ n32490 ;
  assign n32495 = n32335 & ~n32494 ;
  assign n32496 = n32495 ^ n30432 ;
  assign n32497 = n32496 ^ n30428 ;
  assign n32499 = ~n31354 & ~n32498 ;
  assign n32500 = n32499 ^ n31859 ;
  assign n32501 = n32500 ^ n32496 ;
  assign n32502 = ~n32497 & n32501 ;
  assign n32503 = n32502 ^ n30428 ;
  assign n32699 = n32503 ^ n32329 ;
  assign n32700 = ~n32330 & ~n32699 ;
  assign n32701 = n32700 ^ n30404 ;
  assign n32756 = n32710 ^ n32701 ;
  assign n32764 = n32763 ^ n32762 ;
  assign n32765 = ~n31413 & n32764 ;
  assign n32766 = n32765 ^ n31934 ;
  assign n32767 = n32766 ^ n30573 ;
  assign n32768 = n32767 ^ n32766 ;
  assign n32769 = n32768 ^ n32710 ;
  assign n32770 = ~n32756 & n32769 ;
  assign n32771 = n32770 ^ n32767 ;
  assign n32783 = n32766 ^ n30580 ;
  assign n32784 = ~n32771 & ~n32783 ;
  assign n32785 = n32784 ^ n30580 ;
  assign n32882 = n32794 ^ n32785 ;
  assign n32883 = n32795 & n32882 ;
  assign n32884 = n32883 ^ n30424 ;
  assign n32878 = n32877 ^ n32874 ;
  assign n32879 = n31456 & n32878 ;
  assign n32880 = n32879 ^ n32035 ;
  assign n32964 = n32884 ^ n32880 ;
  assign n32972 = n32971 ^ n32970 ;
  assign n32973 = ~n31483 & ~n32972 ;
  assign n32974 = n32973 ^ n31926 ;
  assign n32975 = n32974 ^ n30601 ;
  assign n32976 = n32975 ^ n32884 ;
  assign n32977 = n32976 ^ n32974 ;
  assign n32978 = ~n32964 & ~n32977 ;
  assign n32979 = n32978 ^ n32975 ;
  assign n33024 = n32974 ^ n30611 ;
  assign n33025 = n32979 & ~n33024 ;
  assign n33026 = n33025 ^ n30611 ;
  assign n33073 = n33035 ^ n33026 ;
  assign n33074 = n33035 ^ n30624 ;
  assign n33075 = ~n33073 & n33074 ;
  assign n33076 = n33075 ^ n30624 ;
  assign n33169 = n33086 ^ n33076 ;
  assign n33170 = n33087 & n33169 ;
  assign n33166 = n32069 ^ n30636 ;
  assign n33167 = n33166 ^ n30646 ;
  assign n33168 = n33167 ^ x472 ;
  assign n33171 = n33170 ^ n33168 ;
  assign n33161 = n32214 ^ n32212 ;
  assign n33162 = n33161 ^ n32069 ;
  assign n33163 = n33162 ^ n33083 ;
  assign n33159 = n33083 ^ n32054 ;
  assign n33160 = n33082 & n33159 ;
  assign n33164 = n33163 ^ n33160 ;
  assign n33165 = n31571 & n33164 ;
  assign n33172 = n33171 ^ n33165 ;
  assign n32980 = n32979 ^ n30611 ;
  assign n32981 = n32980 ^ x475 ;
  assign n32881 = n32880 ^ n30601 ;
  assign n32885 = n32884 ^ n32881 ;
  assign n32886 = n32885 ^ x476 ;
  assign n32796 = n32795 ^ n32785 ;
  assign n32797 = n32796 ^ x477 ;
  assign n32772 = n32771 ^ n30580 ;
  assign n32773 = n32772 ^ x478 ;
  assign n32702 = n32701 ^ n30573 ;
  assign n32711 = n32710 ^ n32702 ;
  assign n32712 = n32711 ^ x479 ;
  assign n32504 = n32503 ^ n32330 ;
  assign n32505 = n32504 ^ x464 ;
  assign n32506 = n32500 ^ n32497 ;
  assign n32507 = n32506 ^ x465 ;
  assign n32508 = n32485 ^ n30435 ;
  assign n32509 = n32508 ^ n32488 ;
  assign n32510 = n32509 ^ x467 ;
  assign n32622 = n32621 ^ n32511 ;
  assign n32623 = n32621 ^ x468 ;
  assign n32624 = n32622 & n32623 ;
  assign n32625 = n32624 ^ x468 ;
  assign n32626 = n32625 ^ n32509 ;
  assign n32627 = ~n32510 & n32626 ;
  assign n32628 = n32627 ^ x467 ;
  assign n32629 = n32628 ^ x466 ;
  assign n32630 = n32494 ^ n30432 ;
  assign n32631 = n32630 ^ n32628 ;
  assign n32632 = n32629 & ~n32631 ;
  assign n32633 = n32632 ^ x466 ;
  assign n32634 = n32633 ^ n32506 ;
  assign n32635 = n32507 & ~n32634 ;
  assign n32636 = n32635 ^ x465 ;
  assign n32696 = n32636 ^ n32504 ;
  assign n32697 = n32505 & ~n32696 ;
  assign n32698 = n32697 ^ x464 ;
  assign n32753 = n32711 ^ n32698 ;
  assign n32754 = n32712 & ~n32753 ;
  assign n32755 = n32754 ^ x479 ;
  assign n32780 = n32772 ^ n32755 ;
  assign n32781 = ~n32773 & n32780 ;
  assign n32782 = n32781 ^ x478 ;
  assign n32887 = n32796 ^ n32782 ;
  assign n32888 = ~n32797 & n32887 ;
  assign n32889 = n32888 ^ x477 ;
  assign n32961 = n32889 ^ n32885 ;
  assign n32962 = ~n32886 & n32961 ;
  assign n32963 = n32962 ^ x476 ;
  assign n33038 = n32980 ^ n32963 ;
  assign n33039 = n32981 & ~n33038 ;
  assign n33040 = n33039 ^ x475 ;
  assign n33027 = n33026 ^ n30624 ;
  assign n33036 = n33035 ^ n33027 ;
  assign n33072 = n33040 ^ n33036 ;
  assign n33088 = n33087 ^ n33076 ;
  assign n33089 = n33088 ^ x474 ;
  assign n33090 = n33089 ^ n33036 ;
  assign n33091 = n33090 ^ n33088 ;
  assign n33092 = n33072 & ~n33091 ;
  assign n33093 = n33092 ^ n33089 ;
  assign n32637 = n32636 ^ n32505 ;
  assign n32638 = n32633 ^ n32507 ;
  assign n32639 = n32630 ^ n32629 ;
  assign n32640 = n32625 ^ n32510 ;
  assign n32691 = ~n32688 & ~n32690 ;
  assign n32692 = n32640 & ~n32691 ;
  assign n32693 = n32639 & ~n32692 ;
  assign n32694 = n32638 & n32693 ;
  assign n32695 = ~n32637 & ~n32694 ;
  assign n32713 = n32712 ^ n32698 ;
  assign n32752 = n32695 & ~n32713 ;
  assign n32774 = n32773 ^ n32755 ;
  assign n32779 = n32752 & n32774 ;
  assign n32798 = n32797 ^ n32782 ;
  assign n32872 = ~n32779 & ~n32798 ;
  assign n32890 = n32889 ^ n32886 ;
  assign n32960 = ~n32872 & n32890 ;
  assign n32982 = n32981 ^ n32963 ;
  assign n33023 = ~n32960 & n32982 ;
  assign n33037 = n33036 ^ x474 ;
  assign n33041 = n33040 ^ n33037 ;
  assign n33095 = ~n33023 & n33041 ;
  assign n33154 = n33095 ^ n33088 ;
  assign n33157 = n33093 & ~n33154 ;
  assign n33153 = n33093 ^ n33088 ;
  assign n33155 = n33154 ^ n33153 ;
  assign n33156 = ~x473 & n33155 ;
  assign n33158 = n33157 ^ n33156 ;
  assign n33173 = n33172 ^ n33158 ;
  assign n33174 = n33173 ^ n32349 ;
  assign n32983 = n32982 ^ n32960 ;
  assign n32984 = n32983 ^ n32358 ;
  assign n32891 = n32890 ^ n32872 ;
  assign n32892 = n32891 ^ n32436 ;
  assign n32799 = n32798 ^ n32779 ;
  assign n32800 = n32799 ^ n32362 ;
  assign n32714 = n32713 ^ n32695 ;
  assign n32715 = n32714 ^ n32369 ;
  assign n32716 = n32691 ^ n32640 ;
  assign n32717 = n32716 ^ n32385 ;
  assign n32726 = n32725 ^ n32718 ;
  assign n32727 = n32725 ^ n32403 ;
  assign n32728 = ~n32726 & n32727 ;
  assign n32729 = n32728 ^ n32403 ;
  assign n32730 = n32729 ^ n32716 ;
  assign n32731 = ~n32717 & ~n32730 ;
  assign n32732 = n32731 ^ n32385 ;
  assign n32733 = n32732 ^ n32382 ;
  assign n32734 = n32692 ^ n32639 ;
  assign n32735 = n32734 ^ n32732 ;
  assign n32736 = n32733 & ~n32735 ;
  assign n32737 = n32736 ^ n32382 ;
  assign n32738 = n32737 ^ n32377 ;
  assign n32739 = n32693 ^ n32638 ;
  assign n32740 = n32739 ^ n32737 ;
  assign n32741 = n32738 & n32740 ;
  assign n32742 = n32741 ^ n32377 ;
  assign n32743 = n32742 ^ n32374 ;
  assign n32744 = n32694 ^ n32637 ;
  assign n32745 = n32744 ^ n32742 ;
  assign n32746 = n32743 & ~n32745 ;
  assign n32747 = n32746 ^ n32374 ;
  assign n32748 = n32747 ^ n32714 ;
  assign n32749 = n32715 & n32748 ;
  assign n32750 = n32749 ^ n32369 ;
  assign n32751 = n32750 ^ n32366 ;
  assign n32775 = n32774 ^ n32752 ;
  assign n32776 = n32775 ^ n32750 ;
  assign n32777 = n32751 & n32776 ;
  assign n32778 = n32777 ^ n32366 ;
  assign n32893 = n32799 ^ n32778 ;
  assign n32894 = n32800 & ~n32893 ;
  assign n32895 = n32894 ^ n32362 ;
  assign n32957 = n32895 ^ n32891 ;
  assign n32958 = n32892 & ~n32957 ;
  assign n32959 = n32958 ^ n32436 ;
  assign n33043 = n32983 ^ n32959 ;
  assign n33044 = ~n32984 & n33043 ;
  assign n33045 = n33044 ^ n32358 ;
  assign n33046 = n33045 ^ n32353 ;
  assign n33042 = n33041 ^ n33023 ;
  assign n33097 = n33045 ^ n33042 ;
  assign n33098 = ~n33046 & ~n33097 ;
  assign n33099 = n33098 ^ n32353 ;
  assign n33100 = n33099 ^ n32450 ;
  assign n33094 = n33093 ^ x473 ;
  assign n33096 = n33095 ^ n33094 ;
  assign n33150 = n33099 ^ n33096 ;
  assign n33151 = n33100 & n33150 ;
  assign n33152 = n33151 ^ n32450 ;
  assign n33204 = n33173 ^ n33152 ;
  assign n33205 = n33174 & ~n33204 ;
  assign n33206 = n33205 ^ n32349 ;
  assign n33207 = n33206 ^ n32346 ;
  assign n33208 = n32643 ^ n32641 ;
  assign n33210 = n33208 ^ n32643 ;
  assign n33211 = n33210 ^ n33206 ;
  assign n33212 = n33207 & ~n33211 ;
  assign n33213 = n33212 ^ n32643 ;
  assign n33240 = n32646 ^ n32644 ;
  assign n33242 = n33240 ^ n32465 ;
  assign n33241 = n33240 ^ n33208 ;
  assign n33243 = n33242 ^ n33241 ;
  assign n33244 = n33213 & ~n33243 ;
  assign n33245 = n33244 ^ n33242 ;
  assign n33292 = n32475 ^ n32341 ;
  assign n33291 = n33240 ^ n32475 ;
  assign n33293 = n33292 ^ n33291 ;
  assign n33294 = n33245 & ~n33293 ;
  assign n33295 = n33294 ^ n33292 ;
  assign n33311 = n32475 ^ n32336 ;
  assign n33296 = n32649 ^ n32647 ;
  assign n33310 = n33296 ^ n32336 ;
  assign n33312 = n33311 ^ n33310 ;
  assign n33313 = ~n33295 & ~n33312 ;
  assign n33314 = n33313 ^ n33311 ;
  assign n33315 = n32651 ^ n32650 ;
  assign n33354 = n33315 ^ n32336 ;
  assign n33355 = ~n33314 & ~n33354 ;
  assign n33356 = n33355 ^ n32336 ;
  assign n33357 = n33356 ^ n32486 ;
  assign n33358 = ~n33353 & n33357 ;
  assign n33359 = n33358 ^ n33352 ;
  assign n33360 = n33359 ^ n32332 ;
  assign n33361 = ~n33351 & n33360 ;
  assign n33362 = n33361 ^ n33350 ;
  assign n33364 = n33363 ^ n33362 ;
  assign n33365 = n33363 ^ n32498 ;
  assign n33366 = n33364 & ~n33365 ;
  assign n33368 = n33367 ^ n33366 ;
  assign n33399 = n33369 ^ n33368 ;
  assign n33401 = n33400 ^ n33399 ;
  assign n33411 = n33365 ^ n33362 ;
  assign n33665 = n33411 ^ n33399 ;
  assign n33473 = n32677 ^ n32675 ;
  assign n33474 = n33473 ^ n33033 ;
  assign n33460 = n32674 ^ n32673 ;
  assign n33461 = n33460 ^ n32972 ;
  assign n33385 = n32672 ^ n32670 ;
  assign n33386 = n33385 ^ n32878 ;
  assign n33346 = n32669 ^ n32667 ;
  assign n33347 = n33346 ^ n32792 ;
  assign n33348 = n32666 ^ n32664 ;
  assign n33349 = n33348 ^ n32764 ;
  assign n33373 = n32663 ^ n32662 ;
  assign n33370 = n33369 ^ n32327 ;
  assign n33371 = n33368 & ~n33370 ;
  assign n33372 = n33371 ^ n32327 ;
  assign n33374 = n33373 ^ n33372 ;
  assign n33375 = n33348 ^ n32708 ;
  assign n33376 = n33375 ^ n33372 ;
  assign n33377 = n33376 ^ n33348 ;
  assign n33378 = n33374 & ~n33377 ;
  assign n33379 = n33378 ^ n33375 ;
  assign n33380 = n33349 & ~n33379 ;
  assign n33381 = n33380 ^ n32764 ;
  assign n33382 = n33381 ^ n33346 ;
  assign n33383 = n33347 & ~n33382 ;
  assign n33384 = n33383 ^ n32792 ;
  assign n33457 = n33385 ^ n33384 ;
  assign n33458 = ~n33386 & n33457 ;
  assign n33459 = n33458 ^ n32878 ;
  assign n33470 = n33460 ^ n33459 ;
  assign n33471 = n33461 & n33470 ;
  assign n33472 = n33471 ^ n32972 ;
  assign n33539 = n33473 ^ n33472 ;
  assign n33540 = ~n33474 & n33539 ;
  assign n33541 = n33540 ^ n33033 ;
  assign n33537 = n32679 ^ n32678 ;
  assign n33538 = n33537 ^ n33084 ;
  assign n33542 = n33541 ^ n33538 ;
  assign n33543 = ~n32054 & n33542 ;
  assign n33544 = n33543 ^ n33084 ;
  assign n33545 = n33544 ^ n31525 ;
  assign n33475 = n33474 ^ n33472 ;
  assign n33476 = n31921 & n33475 ;
  assign n33477 = n33476 ^ n33033 ;
  assign n33533 = n33477 ^ n31503 ;
  assign n33462 = n33461 ^ n33459 ;
  assign n33463 = ~n31926 & n33462 ;
  assign n33464 = n33463 ^ n32972 ;
  assign n33387 = n33386 ^ n33384 ;
  assign n33402 = ~n32035 & ~n33387 ;
  assign n33403 = n33402 ^ n32878 ;
  assign n33404 = n33403 ^ n31456 ;
  assign n33390 = n33381 ^ n33347 ;
  assign n33448 = ~n31931 & n33390 ;
  assign n33449 = n33448 ^ n32792 ;
  assign n33393 = n33379 ^ n32764 ;
  assign n33405 = ~n31934 & n33393 ;
  assign n33406 = n33405 ^ n32764 ;
  assign n33407 = n33406 ^ n31413 ;
  assign n33408 = n31942 & n33399 ;
  assign n33409 = n33408 ^ n32327 ;
  assign n33410 = n33409 ^ n31024 ;
  assign n33412 = n31859 & n33411 ;
  assign n33413 = n33412 ^ n32498 ;
  assign n33414 = n33413 ^ n31354 ;
  assign n33425 = n33359 ^ n33351 ;
  assign n33426 = ~n32008 & n33425 ;
  assign n33427 = n33426 ^ n32332 ;
  assign n33101 = n33100 ^ n33096 ;
  assign n33102 = n31965 & ~n33101 ;
  assign n33103 = n33102 ^ n32450 ;
  assign n33104 = n33103 ^ n31217 ;
  assign n33047 = n33046 ^ n33042 ;
  assign n33048 = n31766 & n33047 ;
  assign n33049 = n33048 ^ n32353 ;
  assign n33050 = n33049 ^ n31200 ;
  assign n32861 = n32775 ^ n32751 ;
  assign n32862 = n31602 & n32861 ;
  assign n32863 = n32862 ^ n32366 ;
  assign n32803 = n32747 ^ n32715 ;
  assign n32804 = n31654 & n32803 ;
  assign n32805 = n32804 ^ n32369 ;
  assign n32806 = n32805 ^ n31118 ;
  assign n32821 = n32820 ^ n32810 ;
  assign n32822 = n32729 ^ n32717 ;
  assign n32823 = n31618 & n32822 ;
  assign n32824 = n32823 ^ n32385 ;
  assign n32825 = n32824 ^ n31049 ;
  assign n32826 = n32825 ^ n32810 ;
  assign n32827 = n32826 ^ n32824 ;
  assign n32828 = ~n32821 & n32827 ;
  assign n32829 = n32828 ^ n32825 ;
  assign n32830 = n32734 ^ n32733 ;
  assign n32831 = n31614 & n32830 ;
  assign n32832 = n32831 ^ n32382 ;
  assign n32834 = n32832 ^ n31060 ;
  assign n32833 = n32832 ^ n32824 ;
  assign n32835 = n32834 ^ n32833 ;
  assign n32836 = n32829 & ~n32835 ;
  assign n32837 = n32836 ^ n32834 ;
  assign n32838 = n32739 ^ n32738 ;
  assign n32839 = n31610 & ~n32838 ;
  assign n32840 = n32839 ^ n32377 ;
  assign n32842 = n32840 ^ n31071 ;
  assign n32841 = n32840 ^ n32832 ;
  assign n32843 = n32842 ^ n32841 ;
  assign n32844 = n32837 & ~n32843 ;
  assign n32845 = n32844 ^ n32842 ;
  assign n32846 = n32744 ^ n32743 ;
  assign n32847 = n31606 & n32846 ;
  assign n32848 = n32847 ^ n32374 ;
  assign n32850 = n32848 ^ n31088 ;
  assign n32849 = n32848 ^ n32840 ;
  assign n32851 = n32850 ^ n32849 ;
  assign n32852 = n32845 & n32851 ;
  assign n32853 = n32852 ^ n32850 ;
  assign n32855 = n32805 ^ n31030 ;
  assign n32854 = n32848 ^ n32805 ;
  assign n32856 = n32855 ^ n32854 ;
  assign n32857 = ~n32853 & ~n32856 ;
  assign n32858 = n32857 ^ n32855 ;
  assign n32859 = n32806 & ~n32858 ;
  assign n32860 = n32859 ^ n31118 ;
  assign n32864 = n32863 ^ n32860 ;
  assign n32801 = n32800 ^ n32778 ;
  assign n32865 = ~n31599 & ~n32801 ;
  assign n32866 = n32865 ^ n32362 ;
  assign n32867 = n32866 ^ n31136 ;
  assign n32868 = n32867 ^ n32860 ;
  assign n32869 = n32868 ^ n32866 ;
  assign n32870 = ~n32864 & ~n32869 ;
  assign n32871 = n32870 ^ n32867 ;
  assign n32896 = n32895 ^ n32892 ;
  assign n32897 = ~n31672 & ~n32896 ;
  assign n32898 = n32897 ^ n32436 ;
  assign n32900 = n32898 ^ n31151 ;
  assign n32899 = n32898 ^ n32866 ;
  assign n32901 = n32900 ^ n32899 ;
  assign n32902 = n32871 & ~n32901 ;
  assign n32903 = n32902 ^ n32900 ;
  assign n32988 = n32898 ^ n31165 ;
  assign n32989 = n32903 & ~n32988 ;
  assign n32990 = n32989 ^ n31165 ;
  assign n32991 = n32990 ^ n31185 ;
  assign n32985 = n32984 ^ n32959 ;
  assign n32986 = n31745 & n32985 ;
  assign n32987 = n32986 ^ n32358 ;
  assign n33020 = n32990 ^ n32987 ;
  assign n33021 = ~n32991 & n33020 ;
  assign n33022 = n33021 ^ n31185 ;
  assign n33069 = n33049 ^ n33022 ;
  assign n33070 = n33050 & n33069 ;
  assign n33071 = n33070 ^ n31200 ;
  assign n33178 = n33103 ^ n33071 ;
  assign n33179 = n33104 & ~n33178 ;
  assign n33180 = n33179 ^ n31217 ;
  assign n33181 = n33180 ^ n31232 ;
  assign n33175 = n33174 ^ n33152 ;
  assign n33176 = ~n31876 & n33175 ;
  assign n33177 = n33176 ^ n32349 ;
  assign n33218 = n33180 ^ n33177 ;
  assign n33219 = ~n33181 & ~n33218 ;
  assign n33220 = n33219 ^ n31232 ;
  assign n33221 = n33220 ^ n31246 ;
  assign n33222 = n32641 ^ n32346 ;
  assign n33223 = n33222 ^ n33206 ;
  assign n33224 = ~n31957 & n33223 ;
  assign n33225 = n33224 ^ n32346 ;
  assign n33226 = n33225 ^ n33220 ;
  assign n33227 = n33221 & ~n33226 ;
  assign n33228 = n33227 ^ n31246 ;
  assign n33214 = n33213 ^ n32465 ;
  assign n33215 = n31872 & n33214 ;
  assign n33216 = n33215 ^ n32465 ;
  assign n33239 = n33228 ^ n33216 ;
  assign n33246 = n33245 ^ n32341 ;
  assign n33247 = ~n31986 & n33246 ;
  assign n33248 = n33247 ^ n32341 ;
  assign n33249 = n33248 ^ n31262 ;
  assign n33250 = n33249 ^ n33248 ;
  assign n33251 = n33250 ^ n33216 ;
  assign n33252 = ~n33239 & n33251 ;
  assign n33253 = n33252 ^ n33249 ;
  assign n33300 = n33248 ^ n31282 ;
  assign n33301 = ~n33253 & ~n33300 ;
  assign n33302 = n33301 ^ n31282 ;
  assign n33303 = n33302 ^ n31293 ;
  assign n33297 = n33296 ^ n33295 ;
  assign n33298 = n31949 & n33297 ;
  assign n33299 = n33298 ^ n32475 ;
  assign n33319 = n33302 ^ n33299 ;
  assign n33320 = n33303 & ~n33319 ;
  assign n33321 = n33320 ^ n31293 ;
  assign n33322 = n33321 ^ n31312 ;
  assign n33316 = n33315 ^ n33314 ;
  assign n33317 = n31866 & ~n33316 ;
  assign n33318 = n33317 ^ n32336 ;
  assign n33415 = n33321 ^ n33318 ;
  assign n33416 = n33322 & n33415 ;
  assign n33417 = n33416 ^ n31312 ;
  assign n33418 = n33417 ^ n31324 ;
  assign n33419 = n33356 ^ n33353 ;
  assign n33420 = ~n31864 & n33419 ;
  assign n33421 = n33420 ^ n32486 ;
  assign n33422 = n33421 ^ n33417 ;
  assign n33423 = n33418 & ~n33422 ;
  assign n33424 = n33423 ^ n31324 ;
  assign n33428 = n33427 ^ n33424 ;
  assign n33429 = n33413 ^ n31339 ;
  assign n33430 = n33429 ^ n33413 ;
  assign n33431 = n33430 ^ n33424 ;
  assign n33432 = ~n33428 & ~n33431 ;
  assign n33433 = n33432 ^ n33429 ;
  assign n33434 = n33414 & ~n33433 ;
  assign n33435 = n33434 ^ n31354 ;
  assign n33436 = n33435 ^ n33409 ;
  assign n33437 = n33410 & ~n33436 ;
  assign n33438 = n33437 ^ n31024 ;
  assign n33439 = n33438 ^ n31390 ;
  assign n33396 = n33373 ^ n32708 ;
  assign n33397 = n33396 ^ n33372 ;
  assign n33440 = ~n31939 & ~n33397 ;
  assign n33441 = n33440 ^ n32708 ;
  assign n33442 = n33441 ^ n33438 ;
  assign n33443 = n33439 & n33442 ;
  assign n33444 = n33443 ^ n31390 ;
  assign n33445 = n33444 ^ n33406 ;
  assign n33446 = ~n33407 & n33445 ;
  assign n33447 = n33446 ^ n31413 ;
  assign n33450 = n33449 ^ n33447 ;
  assign n33451 = n33449 ^ n31442 ;
  assign n33452 = n33450 & n33451 ;
  assign n33453 = n33452 ^ n31442 ;
  assign n33454 = n33453 ^ n33403 ;
  assign n33455 = n33404 & ~n33454 ;
  assign n33456 = n33455 ^ n31456 ;
  assign n33465 = n33464 ^ n33456 ;
  assign n33466 = n33464 ^ n31483 ;
  assign n33467 = n33465 & n33466 ;
  assign n33468 = n33467 ^ n31483 ;
  assign n33534 = n33477 ^ n33468 ;
  assign n33535 = ~n33533 & ~n33534 ;
  assign n33536 = n33535 ^ n31503 ;
  assign n33546 = n33545 ^ n33536 ;
  assign n33591 = n33546 ^ x185 ;
  assign n33469 = n33468 ^ n31503 ;
  assign n33478 = n33477 ^ n33469 ;
  assign n33479 = n33478 ^ x186 ;
  assign n33525 = n33466 ^ n33456 ;
  assign n33480 = n33453 ^ n33404 ;
  assign n33481 = n33480 ^ x188 ;
  assign n33517 = n33451 ^ n33447 ;
  assign n33482 = n33441 ^ n33439 ;
  assign n33483 = n33482 ^ x191 ;
  assign n33484 = n33433 ^ n31354 ;
  assign n33485 = n33484 ^ x177 ;
  assign n33494 = n33427 ^ n31339 ;
  assign n33495 = n33494 ^ n33424 ;
  assign n33304 = n33303 ^ n33299 ;
  assign n33305 = n33304 ^ x181 ;
  assign n33233 = n33225 ^ n33221 ;
  assign n33182 = n33181 ^ n33177 ;
  assign n33183 = n33182 ^ x169 ;
  assign n32992 = n32991 ^ n32987 ;
  assign n32993 = n32992 ^ x172 ;
  assign n32904 = n32903 ^ n31165 ;
  assign n32905 = n32904 ^ x173 ;
  assign n32949 = n32871 ^ n31151 ;
  assign n32906 = n32860 ^ n31136 ;
  assign n32907 = n32906 ^ n32863 ;
  assign n32908 = n32907 ^ x175 ;
  assign n32909 = n32853 ^ n31030 ;
  assign n32910 = n32909 ^ x161 ;
  assign n32933 = n32845 ^ n31088 ;
  assign n32911 = n32837 ^ n31071 ;
  assign n32912 = n32911 ^ x163 ;
  assign n32925 = n32829 ^ n31060 ;
  assign n32921 = n32920 ^ n32914 ;
  assign n32922 = n32920 ^ x165 ;
  assign n32923 = n32921 & n32922 ;
  assign n32924 = n32923 ^ x165 ;
  assign n32926 = n32925 ^ n32924 ;
  assign n32927 = n32925 ^ x164 ;
  assign n32928 = ~n32926 & n32927 ;
  assign n32929 = n32928 ^ x164 ;
  assign n32930 = n32929 ^ n32911 ;
  assign n32931 = n32912 & ~n32930 ;
  assign n32932 = n32931 ^ x163 ;
  assign n32934 = n32933 ^ n32932 ;
  assign n32935 = n32933 ^ x162 ;
  assign n32936 = n32934 & ~n32935 ;
  assign n32937 = n32936 ^ x162 ;
  assign n32938 = n32937 ^ n32909 ;
  assign n32939 = ~n32910 & n32938 ;
  assign n32940 = n32939 ^ x161 ;
  assign n32941 = n32940 ^ x160 ;
  assign n32942 = n32858 ^ n31118 ;
  assign n32943 = n32942 ^ n32940 ;
  assign n32944 = n32941 & n32943 ;
  assign n32945 = n32944 ^ x160 ;
  assign n32946 = n32945 ^ n32907 ;
  assign n32947 = n32908 & ~n32946 ;
  assign n32948 = n32947 ^ x175 ;
  assign n32950 = n32949 ^ n32948 ;
  assign n32951 = n32949 ^ x174 ;
  assign n32952 = n32950 & ~n32951 ;
  assign n32953 = n32952 ^ x174 ;
  assign n32954 = n32953 ^ n32904 ;
  assign n32955 = ~n32905 & n32954 ;
  assign n32956 = n32955 ^ x173 ;
  assign n33053 = n32992 ^ n32956 ;
  assign n33054 = n32993 & ~n33053 ;
  assign n33055 = n33054 ^ x172 ;
  assign n33051 = n33050 ^ n33022 ;
  assign n33068 = n33055 ^ n33051 ;
  assign n33105 = n33104 ^ n33071 ;
  assign n33106 = n33105 ^ x171 ;
  assign n33107 = n33106 ^ n33105 ;
  assign n33108 = n33107 ^ n33055 ;
  assign n33109 = n33068 & n33108 ;
  assign n33110 = n33109 ^ n33106 ;
  assign n33147 = n33105 ^ x170 ;
  assign n33148 = ~n33110 & n33147 ;
  assign n33149 = n33148 ^ x170 ;
  assign n33230 = n33182 ^ n33149 ;
  assign n33231 = ~n33183 & n33230 ;
  assign n33232 = n33231 ^ x169 ;
  assign n33234 = n33233 ^ n33232 ;
  assign n33235 = n33233 ^ x168 ;
  assign n33236 = n33234 & ~n33235 ;
  assign n33237 = n33236 ^ x168 ;
  assign n33217 = n33216 ^ n31262 ;
  assign n33229 = n33228 ^ n33217 ;
  assign n33238 = n33237 ^ n33229 ;
  assign n33254 = n33253 ^ n31282 ;
  assign n33255 = n33254 ^ x183 ;
  assign n33256 = n33255 ^ n33254 ;
  assign n33257 = n33256 ^ n33229 ;
  assign n33258 = n33238 & ~n33257 ;
  assign n33259 = n33258 ^ n33255 ;
  assign n33288 = n33254 ^ x182 ;
  assign n33289 = ~n33259 & n33288 ;
  assign n33290 = n33289 ^ x182 ;
  assign n33324 = n33304 ^ n33290 ;
  assign n33325 = n33305 & ~n33324 ;
  assign n33326 = n33325 ^ x181 ;
  assign n33327 = n33326 ^ x180 ;
  assign n33323 = n33322 ^ n33318 ;
  assign n33486 = n33326 ^ n33323 ;
  assign n33487 = n33327 & n33486 ;
  assign n33488 = n33487 ^ x180 ;
  assign n33489 = n33488 ^ x179 ;
  assign n33490 = n33421 ^ n33418 ;
  assign n33491 = n33490 ^ n33488 ;
  assign n33492 = n33489 & ~n33491 ;
  assign n33493 = n33492 ^ x179 ;
  assign n33496 = n33495 ^ n33493 ;
  assign n33497 = n33484 ^ x178 ;
  assign n33498 = n33497 ^ n33484 ;
  assign n33499 = n33498 ^ n33493 ;
  assign n33500 = n33496 & n33499 ;
  assign n33501 = n33500 ^ n33497 ;
  assign n33502 = ~n33485 & n33501 ;
  assign n33503 = n33502 ^ x177 ;
  assign n33504 = n33503 ^ x176 ;
  assign n33505 = n33435 ^ n33410 ;
  assign n33506 = n33505 ^ n33503 ;
  assign n33507 = n33504 & n33506 ;
  assign n33508 = n33507 ^ x176 ;
  assign n33509 = n33508 ^ n33482 ;
  assign n33510 = n33483 & ~n33509 ;
  assign n33511 = n33510 ^ x191 ;
  assign n33512 = n33511 ^ x190 ;
  assign n33513 = n33444 ^ n33407 ;
  assign n33514 = n33513 ^ n33511 ;
  assign n33515 = n33512 & ~n33514 ;
  assign n33516 = n33515 ^ x190 ;
  assign n33518 = n33517 ^ n33516 ;
  assign n33519 = n33517 ^ x189 ;
  assign n33520 = n33518 & ~n33519 ;
  assign n33521 = n33520 ^ x189 ;
  assign n33522 = n33521 ^ n33480 ;
  assign n33523 = n33481 & ~n33522 ;
  assign n33524 = n33523 ^ x188 ;
  assign n33526 = n33525 ^ n33524 ;
  assign n33527 = n33525 ^ x187 ;
  assign n33528 = ~n33526 & n33527 ;
  assign n33529 = n33528 ^ x187 ;
  assign n33530 = n33529 ^ n33478 ;
  assign n33531 = n33479 & ~n33530 ;
  assign n33532 = n33531 ^ x186 ;
  assign n33592 = n33591 ^ n33532 ;
  assign n33328 = n33327 ^ n33323 ;
  assign n33306 = n33305 ^ n33290 ;
  assign n33260 = n33259 ^ x182 ;
  assign n33184 = n33183 ^ n33149 ;
  assign n33111 = n33110 ^ x170 ;
  assign n33052 = n33051 ^ x171 ;
  assign n33056 = n33055 ^ n33052 ;
  assign n32994 = n32993 ^ n32956 ;
  assign n33000 = ~n32996 & n32999 ;
  assign n33001 = n32927 ^ n32924 ;
  assign n33002 = ~n33000 & ~n33001 ;
  assign n33003 = n32929 ^ n32912 ;
  assign n33004 = n33002 & ~n33003 ;
  assign n33005 = n32935 ^ n32932 ;
  assign n33006 = n33004 & n33005 ;
  assign n33007 = n32937 ^ n32910 ;
  assign n33008 = ~n33006 & ~n33007 ;
  assign n33009 = n32942 ^ n32941 ;
  assign n33010 = n33008 & ~n33009 ;
  assign n33011 = n32945 ^ n32908 ;
  assign n33012 = n33010 & n33011 ;
  assign n33013 = n32951 ^ n32948 ;
  assign n33014 = n33012 & ~n33013 ;
  assign n33015 = n32953 ^ n32905 ;
  assign n33016 = n33014 & ~n33015 ;
  assign n33057 = n32994 & n33016 ;
  assign n33112 = ~n33056 & n33057 ;
  assign n33185 = ~n33111 & ~n33112 ;
  assign n33261 = ~n33184 & ~n33185 ;
  assign n33262 = n33235 ^ n33232 ;
  assign n33263 = ~n33261 & n33262 ;
  assign n33264 = n33229 ^ x183 ;
  assign n33265 = n33264 ^ n33237 ;
  assign n33266 = n33263 & n33265 ;
  assign n33307 = ~n33260 & n33266 ;
  assign n33329 = n33306 & ~n33307 ;
  assign n33549 = ~n33328 & n33329 ;
  assign n33550 = n33490 ^ n33489 ;
  assign n33551 = ~n33549 & ~n33550 ;
  assign n33552 = n33495 ^ x178 ;
  assign n33553 = n33552 ^ n33493 ;
  assign n33554 = ~n33551 & ~n33553 ;
  assign n33555 = n33501 ^ x177 ;
  assign n33556 = n33554 & ~n33555 ;
  assign n33557 = n33505 ^ n33504 ;
  assign n33558 = ~n33556 & n33557 ;
  assign n33559 = n33508 ^ n33483 ;
  assign n33560 = ~n33558 & n33559 ;
  assign n33561 = n33513 ^ n33512 ;
  assign n33562 = n33560 & n33561 ;
  assign n33563 = n33519 ^ n33516 ;
  assign n33564 = ~n33562 & n33563 ;
  assign n33565 = n33521 ^ n33481 ;
  assign n33566 = n33564 & ~n33565 ;
  assign n33567 = n33527 ^ n33524 ;
  assign n33568 = n33566 & ~n33567 ;
  assign n33569 = n33529 ^ n33479 ;
  assign n33570 = n33568 & ~n33569 ;
  assign n33593 = n33592 ^ n33570 ;
  assign n33594 = n33593 ^ n33316 ;
  assign n33595 = n33569 ^ n33568 ;
  assign n33596 = n33595 ^ n33297 ;
  assign n33597 = n33567 ^ n33566 ;
  assign n33598 = n33597 ^ n33246 ;
  assign n33637 = n33565 ^ n33564 ;
  assign n33599 = n33563 ^ n33562 ;
  assign n33600 = n33599 ^ n33223 ;
  assign n33601 = n33561 ^ n33560 ;
  assign n33602 = n33601 ^ n33175 ;
  assign n33603 = n33559 ^ n33558 ;
  assign n33604 = n33603 ^ n33101 ;
  assign n33605 = n33557 ^ n33556 ;
  assign n33606 = n33605 ^ n33047 ;
  assign n33607 = n33555 ^ n33554 ;
  assign n33608 = n33607 ^ n32985 ;
  assign n33609 = n33553 ^ n33551 ;
  assign n33610 = n33609 ^ n32896 ;
  assign n33611 = n33550 ^ n33549 ;
  assign n33612 = n33611 ^ n32801 ;
  assign n33308 = n33307 ^ n33306 ;
  assign n33267 = n33266 ^ n33260 ;
  assign n33268 = n33267 ^ n32846 ;
  assign n33279 = n33265 ^ n33263 ;
  assign n33269 = n33262 ^ n33261 ;
  assign n33270 = n33269 ^ n32830 ;
  assign n33058 = n33057 ^ n33056 ;
  assign n33017 = n33016 ^ n32994 ;
  assign n33018 = n32802 & n33017 ;
  assign n33067 = n33058 ^ n33018 ;
  assign n33113 = n33112 ^ n33111 ;
  assign n33114 = n33113 ^ n32815 ;
  assign n33115 = n33114 ^ n33113 ;
  assign n33116 = n33115 ^ n33058 ;
  assign n33117 = n33067 & n33116 ;
  assign n33118 = n33117 ^ n33114 ;
  assign n33188 = n33113 ^ n32808 ;
  assign n33189 = ~n33118 & ~n33188 ;
  assign n33190 = n33189 ^ n32808 ;
  assign n33186 = n33185 ^ n33184 ;
  assign n33271 = n33190 ^ n33186 ;
  assign n33272 = n33269 ^ n32822 ;
  assign n33273 = n33272 ^ n33269 ;
  assign n33274 = n33273 ^ n33186 ;
  assign n33275 = ~n33271 & ~n33274 ;
  assign n33276 = n33275 ^ n33272 ;
  assign n33277 = ~n33270 & n33276 ;
  assign n33278 = n33277 ^ n32830 ;
  assign n33280 = n33279 ^ n33278 ;
  assign n33281 = n33267 ^ n32838 ;
  assign n33282 = n33281 ^ n33267 ;
  assign n33283 = n33282 ^ n33278 ;
  assign n33284 = ~n33280 & ~n33283 ;
  assign n33285 = n33284 ^ n33281 ;
  assign n33286 = ~n33268 & ~n33285 ;
  assign n33287 = n33286 ^ n32846 ;
  assign n33309 = n33308 ^ n33287 ;
  assign n33330 = n33329 ^ n33328 ;
  assign n33331 = n33330 ^ n32803 ;
  assign n33332 = n33331 ^ n33330 ;
  assign n33333 = n33332 ^ n33287 ;
  assign n33334 = ~n33309 & n33333 ;
  assign n33335 = n33334 ^ n33331 ;
  assign n33613 = n33330 ^ n32861 ;
  assign n33614 = ~n33335 & n33613 ;
  assign n33615 = n33614 ^ n32861 ;
  assign n33616 = n33615 ^ n33611 ;
  assign n33617 = ~n33612 & ~n33616 ;
  assign n33618 = n33617 ^ n32801 ;
  assign n33619 = n33618 ^ n33609 ;
  assign n33620 = n33610 & ~n33619 ;
  assign n33621 = n33620 ^ n32896 ;
  assign n33622 = n33621 ^ n33607 ;
  assign n33623 = n33608 & n33622 ;
  assign n33624 = n33623 ^ n32985 ;
  assign n33625 = n33624 ^ n33605 ;
  assign n33626 = ~n33606 & n33625 ;
  assign n33627 = n33626 ^ n33047 ;
  assign n33628 = n33627 ^ n33603 ;
  assign n33629 = ~n33604 & ~n33628 ;
  assign n33630 = n33629 ^ n33101 ;
  assign n33631 = n33630 ^ n33601 ;
  assign n33632 = ~n33602 & ~n33631 ;
  assign n33633 = n33632 ^ n33175 ;
  assign n33634 = n33633 ^ n33599 ;
  assign n33635 = ~n33600 & n33634 ;
  assign n33636 = n33635 ^ n33223 ;
  assign n33638 = n33637 ^ n33636 ;
  assign n33639 = n33597 ^ n33214 ;
  assign n33640 = n33639 ^ n33597 ;
  assign n33641 = n33640 ^ n33636 ;
  assign n33642 = n33638 & n33641 ;
  assign n33643 = n33642 ^ n33639 ;
  assign n33644 = ~n33598 & n33643 ;
  assign n33645 = n33644 ^ n33246 ;
  assign n33646 = n33645 ^ n33595 ;
  assign n33647 = ~n33596 & n33646 ;
  assign n33648 = n33647 ^ n33297 ;
  assign n33649 = n33648 ^ n33593 ;
  assign n33650 = n33594 & n33649 ;
  assign n33651 = n33650 ^ n33316 ;
  assign n33585 = n33164 ^ n31525 ;
  assign n33586 = n33585 ^ n31571 ;
  assign n33587 = n33586 ^ x184 ;
  assign n33583 = n33544 ^ n33536 ;
  assign n33584 = n33545 & n33583 ;
  assign n33588 = n33587 ^ n33584 ;
  assign n33578 = n32682 ^ n32680 ;
  assign n33579 = n33578 ^ n33164 ;
  assign n33580 = n33579 ^ n33084 ;
  assign n33576 = n33541 ^ n33084 ;
  assign n33577 = ~n33538 & n33576 ;
  assign n33581 = n33580 ^ n33577 ;
  assign n33582 = ~n32069 & n33581 ;
  assign n33589 = n33588 ^ n33582 ;
  assign n33547 = n33546 ^ n33532 ;
  assign n33571 = n33570 ^ n33532 ;
  assign n33574 = ~n33547 & n33571 ;
  assign n33572 = n33571 ^ n33546 ;
  assign n33573 = x185 & n33572 ;
  assign n33575 = n33574 ^ n33573 ;
  assign n33590 = n33589 ^ n33575 ;
  assign n33652 = n33651 ^ n33590 ;
  assign n33653 = n33651 ^ n33419 ;
  assign n33654 = n33652 & ~n33653 ;
  assign n33655 = n33654 ^ n33419 ;
  assign n33656 = n33655 ^ n33425 ;
  assign n33657 = n33411 ^ n32997 ;
  assign n33658 = n33657 ^ n33411 ;
  assign n33659 = n33658 ^ n33655 ;
  assign n33660 = ~n33656 & n33659 ;
  assign n33661 = n33660 ^ n33657 ;
  assign n33662 = n32998 ^ n32997 ;
  assign n33663 = n33662 ^ n33411 ;
  assign n33664 = n33661 & ~n33663 ;
  assign n33666 = n33665 ^ n33664 ;
  assign n33667 = n33401 & ~n33666 ;
  assign n33668 = n33667 ^ n33400 ;
  assign n33395 = n33001 ^ n33000 ;
  assign n33398 = n33397 ^ n33395 ;
  assign n33704 = n33668 ^ n33398 ;
  assign n33705 = ~n32708 & ~n33704 ;
  assign n33706 = n33705 ^ n33397 ;
  assign n33707 = n33706 ^ n31939 ;
  assign n33708 = n33666 ^ n33400 ;
  assign n33709 = n32327 & n33708 ;
  assign n33710 = n33709 ^ n33399 ;
  assign n33711 = n33710 ^ n31942 ;
  assign n33712 = n33662 ^ n33661 ;
  assign n33713 = n32498 & ~n33712 ;
  assign n33714 = n33713 ^ n33411 ;
  assign n33715 = n33714 ^ n31859 ;
  assign n33716 = n33425 ^ n32997 ;
  assign n33717 = n33716 ^ n33655 ;
  assign n33718 = ~n32332 & n33717 ;
  assign n33719 = n33718 ^ n33425 ;
  assign n33720 = n33719 ^ n32008 ;
  assign n33721 = n33590 ^ n33419 ;
  assign n33722 = n33721 ^ n33651 ;
  assign n33723 = ~n32486 & ~n33722 ;
  assign n33724 = n33723 ^ n33419 ;
  assign n33725 = n33724 ^ n31864 ;
  assign n33726 = n33648 ^ n33316 ;
  assign n33727 = n33726 ^ n33593 ;
  assign n33728 = n32336 & n33727 ;
  assign n33729 = n33728 ^ n33316 ;
  assign n33730 = n33729 ^ n31866 ;
  assign n33731 = n33645 ^ n33596 ;
  assign n33732 = ~n32475 & ~n33731 ;
  assign n33733 = n33732 ^ n33297 ;
  assign n33734 = n33733 ^ n31949 ;
  assign n33735 = n33643 ^ n33246 ;
  assign n33736 = n32341 & ~n33735 ;
  assign n33737 = n33736 ^ n33246 ;
  assign n33738 = n33737 ^ n31986 ;
  assign n33739 = n33637 ^ n33214 ;
  assign n33740 = n33739 ^ n33636 ;
  assign n33741 = n32465 & ~n33740 ;
  assign n33742 = n33741 ^ n33214 ;
  assign n33743 = n33742 ^ n31872 ;
  assign n33744 = n33633 ^ n33600 ;
  assign n33745 = n32346 & ~n33744 ;
  assign n33746 = n33745 ^ n33223 ;
  assign n33747 = n33746 ^ n31957 ;
  assign n33823 = n33630 ^ n33602 ;
  assign n33824 = ~n32349 & n33823 ;
  assign n33825 = n33824 ^ n33175 ;
  assign n33752 = n33624 ^ n33606 ;
  assign n33753 = ~n32353 & ~n33752 ;
  assign n33754 = n33753 ^ n33047 ;
  assign n33755 = n33754 ^ n31766 ;
  assign n33756 = n33621 ^ n33608 ;
  assign n33757 = n32358 & ~n33756 ;
  assign n33758 = n33757 ^ n32985 ;
  assign n33759 = n33758 ^ n31745 ;
  assign n33805 = n33618 ^ n33610 ;
  assign n33806 = n32436 & ~n33805 ;
  assign n33807 = n33806 ^ n32896 ;
  assign n33760 = n33615 ^ n33612 ;
  assign n33761 = n32362 & ~n33760 ;
  assign n33762 = n33761 ^ n32801 ;
  assign n33763 = n33762 ^ n31599 ;
  assign n33338 = n33308 ^ n32803 ;
  assign n33339 = n33338 ^ n33287 ;
  assign n33766 = n32369 & n33339 ;
  assign n33767 = n33766 ^ n32803 ;
  assign n33768 = n33767 ^ n31654 ;
  assign n33342 = n33285 ^ n32846 ;
  assign n33769 = ~n32374 & n33342 ;
  assign n33770 = n33769 ^ n32846 ;
  assign n33771 = n33770 ^ n31606 ;
  assign n33783 = n33279 ^ n32838 ;
  assign n33784 = n33783 ^ n33278 ;
  assign n33785 = ~n32377 & ~n33784 ;
  assign n33786 = n33785 ^ n32838 ;
  assign n33772 = n33276 ^ n32830 ;
  assign n33773 = ~n32382 & ~n33772 ;
  assign n33774 = n33773 ^ n32830 ;
  assign n33775 = n33774 ^ n31614 ;
  assign n33062 = n33017 ^ n32802 ;
  assign n33063 = n32390 & ~n33062 ;
  assign n33064 = n33063 ^ n32802 ;
  assign n33065 = n31628 & ~n33064 ;
  assign n33019 = n33018 ^ n32815 ;
  assign n33059 = n33058 ^ n33019 ;
  assign n33060 = n32395 & ~n33059 ;
  assign n33061 = n33060 ^ n32815 ;
  assign n33066 = n33065 ^ n33061 ;
  assign n33119 = n33118 ^ n32808 ;
  assign n33120 = n32403 & ~n33119 ;
  assign n33121 = n33120 ^ n32808 ;
  assign n33122 = n33121 ^ n31625 ;
  assign n33123 = n33122 ^ n33121 ;
  assign n33124 = n33123 ^ n33061 ;
  assign n33125 = ~n33066 & n33124 ;
  assign n33126 = n33125 ^ n33122 ;
  assign n33195 = n33121 ^ n31622 ;
  assign n33196 = n33126 & n33195 ;
  assign n33197 = n33196 ^ n31622 ;
  assign n33187 = n33186 ^ n32822 ;
  assign n33191 = n33190 ^ n33187 ;
  assign n33192 = ~n32385 & n33191 ;
  assign n33193 = n33192 ^ n32822 ;
  assign n33776 = n33197 ^ n33193 ;
  assign n33777 = n33197 ^ n31618 ;
  assign n33778 = n33776 & ~n33777 ;
  assign n33779 = n33778 ^ n31618 ;
  assign n33780 = n33779 ^ n33774 ;
  assign n33781 = n33775 & ~n33780 ;
  assign n33782 = n33781 ^ n31614 ;
  assign n33787 = n33786 ^ n33782 ;
  assign n33788 = n33770 ^ n31610 ;
  assign n33789 = n33788 ^ n33782 ;
  assign n33790 = n33789 ^ n33770 ;
  assign n33791 = n33787 & n33790 ;
  assign n33792 = n33791 ^ n33788 ;
  assign n33793 = n33771 & ~n33792 ;
  assign n33794 = n33793 ^ n31606 ;
  assign n33795 = n33794 ^ n33767 ;
  assign n33796 = n33768 & ~n33795 ;
  assign n33797 = n33796 ^ n31654 ;
  assign n33336 = n33335 ^ n32861 ;
  assign n33764 = n32366 & n33336 ;
  assign n33765 = n33764 ^ n32861 ;
  assign n33798 = n33797 ^ n33765 ;
  assign n33799 = n33797 ^ n31602 ;
  assign n33800 = ~n33798 & n33799 ;
  assign n33801 = n33800 ^ n31602 ;
  assign n33802 = n33801 ^ n33762 ;
  assign n33803 = n33763 & n33802 ;
  assign n33804 = n33803 ^ n31599 ;
  assign n33808 = n33807 ^ n33804 ;
  assign n33809 = n33758 ^ n31672 ;
  assign n33810 = n33809 ^ n33758 ;
  assign n33811 = n33810 ^ n33804 ;
  assign n33812 = ~n33808 & n33811 ;
  assign n33813 = n33812 ^ n33809 ;
  assign n33814 = n33759 & n33813 ;
  assign n33815 = n33814 ^ n31745 ;
  assign n33816 = n33815 ^ n33754 ;
  assign n33817 = n33755 & ~n33816 ;
  assign n33818 = n33817 ^ n31766 ;
  assign n33748 = n33627 ^ n33101 ;
  assign n33749 = n33748 ^ n33603 ;
  assign n33750 = ~n32450 & ~n33749 ;
  assign n33751 = n33750 ^ n33101 ;
  assign n33819 = n33818 ^ n33751 ;
  assign n33820 = n33818 ^ n31965 ;
  assign n33821 = n33819 & n33820 ;
  assign n33822 = n33821 ^ n31965 ;
  assign n33826 = n33825 ^ n33822 ;
  assign n33827 = n33746 ^ n31876 ;
  assign n33828 = n33827 ^ n33746 ;
  assign n33829 = n33828 ^ n33822 ;
  assign n33830 = ~n33826 & ~n33829 ;
  assign n33831 = n33830 ^ n33827 ;
  assign n33832 = ~n33747 & n33831 ;
  assign n33833 = n33832 ^ n31957 ;
  assign n33834 = n33833 ^ n33742 ;
  assign n33835 = n33743 & n33834 ;
  assign n33836 = n33835 ^ n31872 ;
  assign n33837 = n33836 ^ n33737 ;
  assign n33838 = ~n33738 & ~n33837 ;
  assign n33839 = n33838 ^ n31986 ;
  assign n33840 = n33839 ^ n33733 ;
  assign n33841 = n33734 & n33840 ;
  assign n33842 = n33841 ^ n31949 ;
  assign n33843 = n33842 ^ n33729 ;
  assign n33844 = ~n33730 & n33843 ;
  assign n33845 = n33844 ^ n31866 ;
  assign n33846 = n33845 ^ n33724 ;
  assign n33847 = ~n33725 & ~n33846 ;
  assign n33848 = n33847 ^ n31864 ;
  assign n33849 = n33848 ^ n33719 ;
  assign n33850 = ~n33720 & n33849 ;
  assign n33851 = n33850 ^ n32008 ;
  assign n33852 = n33851 ^ n33714 ;
  assign n33853 = n33715 & n33852 ;
  assign n33854 = n33853 ^ n31859 ;
  assign n33855 = n33854 ^ n33710 ;
  assign n33856 = n33711 & ~n33855 ;
  assign n33857 = n33856 ^ n31942 ;
  assign n33858 = n33857 ^ n33706 ;
  assign n33859 = n33707 & n33858 ;
  assign n33860 = n33859 ^ n31939 ;
  assign n34040 = n33860 ^ n31934 ;
  assign n33671 = n33397 ^ n33393 ;
  assign n33669 = n33668 ^ n33395 ;
  assign n33670 = ~n33398 & ~n33669 ;
  assign n33672 = n33671 ^ n33670 ;
  assign n33392 = n33003 ^ n33002 ;
  assign n33700 = n33672 ^ n33392 ;
  assign n33701 = ~n32764 & n33700 ;
  assign n33702 = n33701 ^ n33393 ;
  assign n34041 = n34040 ^ n33702 ;
  assign n33917 = n33857 ^ n31939 ;
  assign n33918 = n33917 ^ n33706 ;
  assign n33919 = n33918 ^ x415 ;
  assign n33920 = n33854 ^ n31942 ;
  assign n33921 = n33920 ^ n33710 ;
  assign n33922 = n33921 ^ x400 ;
  assign n34021 = n33848 ^ n33720 ;
  assign n33923 = n33845 ^ n33725 ;
  assign n33924 = n33923 ^ x403 ;
  assign n34012 = n33842 ^ n33730 ;
  assign n33925 = n33839 ^ n31949 ;
  assign n33926 = n33925 ^ n33733 ;
  assign n33927 = n33926 ^ x405 ;
  assign n33928 = n33836 ^ n31986 ;
  assign n33929 = n33928 ^ n33737 ;
  assign n33930 = n33929 ^ x406 ;
  assign n33931 = n33833 ^ n33743 ;
  assign n33932 = n33931 ^ x407 ;
  assign n33998 = n33831 ^ n31957 ;
  assign n33935 = n33751 ^ n31965 ;
  assign n33936 = n33935 ^ n33818 ;
  assign n33937 = n33936 ^ x394 ;
  assign n33985 = n33815 ^ n33755 ;
  assign n33938 = n33807 ^ n31672 ;
  assign n33939 = n33938 ^ n33804 ;
  assign n33940 = n33939 ^ x397 ;
  assign n33941 = n33801 ^ n33763 ;
  assign n33942 = n33941 ^ x398 ;
  assign n33945 = n33794 ^ n33768 ;
  assign n33946 = n33945 ^ x384 ;
  assign n33947 = n33792 ^ n31606 ;
  assign n33948 = n33947 ^ x385 ;
  assign n33957 = n33786 ^ n31610 ;
  assign n33958 = n33957 ^ n33782 ;
  assign n33194 = n33193 ^ n31618 ;
  assign n33198 = n33197 ^ n33194 ;
  assign n33129 = n32719 ^ n32233 ;
  assign n33130 = n33129 ^ n33063 ;
  assign n33131 = x391 & ~n33130 ;
  assign n33132 = n33131 ^ x390 ;
  assign n33133 = n33065 ^ n31625 ;
  assign n33134 = n33133 ^ n33061 ;
  assign n33135 = n33134 ^ n33131 ;
  assign n33136 = n33132 & ~n33135 ;
  assign n33137 = n33136 ^ x390 ;
  assign n33127 = n33126 ^ n31622 ;
  assign n33143 = n33137 ^ n33127 ;
  assign n33144 = n33137 ^ x389 ;
  assign n33145 = ~n33143 & n33144 ;
  assign n33146 = n33145 ^ x389 ;
  assign n33199 = n33198 ^ n33146 ;
  assign n33950 = n33146 ^ x388 ;
  assign n33951 = n33199 & n33950 ;
  assign n33952 = n33951 ^ x388 ;
  assign n33949 = n33779 ^ n33775 ;
  assign n33953 = n33952 ^ n33949 ;
  assign n33954 = n33952 ^ x387 ;
  assign n33955 = ~n33953 & n33954 ;
  assign n33956 = n33955 ^ x387 ;
  assign n33959 = n33958 ^ n33956 ;
  assign n33960 = n33947 ^ x386 ;
  assign n33961 = n33960 ^ n33947 ;
  assign n33962 = n33961 ^ n33956 ;
  assign n33963 = n33959 & n33962 ;
  assign n33964 = n33963 ^ n33960 ;
  assign n33965 = n33948 & ~n33964 ;
  assign n33966 = n33965 ^ x385 ;
  assign n33967 = n33966 ^ n33945 ;
  assign n33968 = n33946 & ~n33967 ;
  assign n33969 = n33968 ^ x384 ;
  assign n33943 = n33765 ^ n31602 ;
  assign n33944 = n33943 ^ n33797 ;
  assign n33970 = n33969 ^ n33944 ;
  assign n33971 = n33969 ^ x399 ;
  assign n33972 = ~n33970 & n33971 ;
  assign n33973 = n33972 ^ x399 ;
  assign n33974 = n33973 ^ n33941 ;
  assign n33975 = n33942 & ~n33974 ;
  assign n33976 = n33975 ^ x398 ;
  assign n33977 = n33976 ^ n33939 ;
  assign n33978 = ~n33940 & n33977 ;
  assign n33979 = n33978 ^ x397 ;
  assign n33980 = n33979 ^ x396 ;
  assign n33981 = n33813 ^ n31745 ;
  assign n33982 = n33981 ^ n33979 ;
  assign n33983 = n33980 & n33982 ;
  assign n33984 = n33983 ^ x396 ;
  assign n33986 = n33985 ^ n33984 ;
  assign n33987 = n33936 ^ x395 ;
  assign n33988 = n33987 ^ n33936 ;
  assign n33989 = n33988 ^ n33984 ;
  assign n33990 = ~n33986 & n33989 ;
  assign n33991 = n33990 ^ n33987 ;
  assign n33992 = ~n33937 & n33991 ;
  assign n33993 = n33992 ^ x394 ;
  assign n33933 = n33822 ^ n31876 ;
  assign n33934 = n33933 ^ n33825 ;
  assign n33994 = n33993 ^ n33934 ;
  assign n33995 = n33993 ^ x393 ;
  assign n33996 = n33994 & n33995 ;
  assign n33997 = n33996 ^ x393 ;
  assign n33999 = n33998 ^ n33997 ;
  assign n34000 = n33998 ^ x392 ;
  assign n34001 = ~n33999 & n34000 ;
  assign n34002 = n34001 ^ x392 ;
  assign n34003 = n34002 ^ n33931 ;
  assign n34004 = ~n33932 & n34003 ;
  assign n34005 = n34004 ^ x407 ;
  assign n34006 = n34005 ^ n33929 ;
  assign n34007 = ~n33930 & n34006 ;
  assign n34008 = n34007 ^ x406 ;
  assign n34009 = n34008 ^ n33926 ;
  assign n34010 = ~n33927 & n34009 ;
  assign n34011 = n34010 ^ x405 ;
  assign n34013 = n34012 ^ n34011 ;
  assign n34014 = n33923 ^ x404 ;
  assign n34015 = n34014 ^ n33923 ;
  assign n34016 = n34015 ^ n34011 ;
  assign n34017 = n34013 & n34016 ;
  assign n34018 = n34017 ^ n34014 ;
  assign n34019 = ~n33924 & n34018 ;
  assign n34020 = n34019 ^ x403 ;
  assign n34022 = n34021 ^ n34020 ;
  assign n34023 = n33851 ^ n31859 ;
  assign n34024 = n34023 ^ n33714 ;
  assign n34025 = n34024 ^ x402 ;
  assign n34026 = n34025 ^ n34020 ;
  assign n34027 = n34026 ^ n34024 ;
  assign n34028 = ~n34022 & n34027 ;
  assign n34029 = n34028 ^ n34025 ;
  assign n34031 = n33921 ^ x401 ;
  assign n34030 = n34024 ^ n33921 ;
  assign n34032 = n34031 ^ n34030 ;
  assign n34033 = n34029 & ~n34032 ;
  assign n34034 = n34033 ^ n34031 ;
  assign n34035 = n33922 & ~n34034 ;
  assign n34036 = n34035 ^ x400 ;
  assign n34037 = n34036 ^ n33918 ;
  assign n34038 = n33919 & ~n34037 ;
  assign n34039 = n34038 ^ x415 ;
  assign n34042 = n34041 ^ n34039 ;
  assign n33703 = n33702 ^ n31934 ;
  assign n33861 = n33860 ^ n33702 ;
  assign n33862 = ~n33703 & n33861 ;
  assign n33863 = n33862 ^ n31934 ;
  assign n33394 = n33393 ^ n33392 ;
  assign n33673 = ~n33394 & ~n33672 ;
  assign n33674 = n33673 ^ n33393 ;
  assign n33389 = n33005 ^ n33004 ;
  assign n33391 = n33390 ^ n33389 ;
  assign n33696 = n33674 ^ n33391 ;
  assign n33697 = ~n32792 & n33696 ;
  assign n33698 = n33697 ^ n33390 ;
  assign n33699 = n33698 ^ n31931 ;
  assign n33915 = n33863 ^ n33699 ;
  assign n34043 = n33915 ^ x414 ;
  assign n34044 = n34043 ^ n33915 ;
  assign n34045 = n34044 ^ n34039 ;
  assign n34046 = ~n34042 & n34045 ;
  assign n34047 = n34046 ^ n34043 ;
  assign n34121 = n34047 ^ x413 ;
  assign n34066 = n33997 ^ x392 ;
  assign n34067 = n34066 ^ n33998 ;
  assign n34068 = n33958 ^ x386 ;
  assign n34069 = n34068 ^ n33956 ;
  assign n33200 = n33199 ^ x388 ;
  assign n33128 = n33127 ^ x389 ;
  assign n33138 = n33137 ^ n33128 ;
  assign n33139 = n33130 ^ x391 ;
  assign n33140 = n33134 ^ n33132 ;
  assign n33141 = n33139 & ~n33140 ;
  assign n33201 = n33138 & ~n33141 ;
  assign n34070 = ~n33200 & n33201 ;
  assign n34071 = n33949 ^ x387 ;
  assign n34072 = n34071 ^ n33952 ;
  assign n34073 = n34070 & n34072 ;
  assign n34074 = ~n34069 & n34073 ;
  assign n34075 = n33964 ^ x385 ;
  assign n34076 = ~n34074 & ~n34075 ;
  assign n34077 = n33966 ^ n33946 ;
  assign n34078 = n34076 & ~n34077 ;
  assign n34079 = n33944 ^ x399 ;
  assign n34080 = n34079 ^ n33969 ;
  assign n34081 = n34078 & ~n34080 ;
  assign n34082 = n33973 ^ n33942 ;
  assign n34083 = ~n34081 & n34082 ;
  assign n34084 = n33976 ^ n33940 ;
  assign n34085 = n34083 & ~n34084 ;
  assign n34086 = n33981 ^ n33980 ;
  assign n34087 = ~n34085 & n34086 ;
  assign n34088 = n33984 ^ x395 ;
  assign n34089 = n34088 ^ n33985 ;
  assign n34090 = n34087 & ~n34089 ;
  assign n34091 = n33991 ^ x394 ;
  assign n34092 = ~n34090 & ~n34091 ;
  assign n34093 = n33934 ^ x393 ;
  assign n34094 = n34093 ^ n33993 ;
  assign n34095 = ~n34092 & n34094 ;
  assign n34096 = n34067 & ~n34095 ;
  assign n34097 = n34002 ^ x407 ;
  assign n34098 = n34097 ^ n33931 ;
  assign n34099 = ~n34096 & n34098 ;
  assign n34100 = n34005 ^ n33930 ;
  assign n34101 = n34099 & n34100 ;
  assign n34102 = n34008 ^ n33927 ;
  assign n34103 = ~n34101 & ~n34102 ;
  assign n34104 = n34011 ^ x404 ;
  assign n34105 = n34104 ^ n34012 ;
  assign n34106 = ~n34103 & n34105 ;
  assign n34107 = n34018 ^ x403 ;
  assign n34108 = n34106 & n34107 ;
  assign n34109 = n34021 ^ x402 ;
  assign n34110 = n34109 ^ n34020 ;
  assign n34111 = ~n34108 & n34110 ;
  assign n34112 = n34029 ^ x401 ;
  assign n34113 = ~n34111 & n34112 ;
  assign n34114 = n34034 ^ x400 ;
  assign n34115 = ~n34113 & n34114 ;
  assign n34116 = n34036 ^ n33919 ;
  assign n34117 = ~n34115 & ~n34116 ;
  assign n34118 = n34041 ^ x414 ;
  assign n34119 = n34118 ^ n34039 ;
  assign n34120 = ~n34117 & n34119 ;
  assign n34135 = n34121 ^ n34120 ;
  assign n34188 = n34135 ^ n33062 ;
  assign n34258 = n33017 ^ n32719 ;
  assign n34189 = n32802 & n34188 ;
  assign n34259 = n34258 ^ n34189 ;
  assign n34260 = x103 & ~n34259 ;
  assign n34261 = n34260 ^ x102 ;
  assign n33916 = n33915 ^ x413 ;
  assign n34048 = n33916 & ~n34047 ;
  assign n34049 = n34048 ^ x413 ;
  assign n33864 = n33863 ^ n33698 ;
  assign n33865 = ~n33699 & n33864 ;
  assign n33866 = n33865 ^ n31931 ;
  assign n33912 = n33866 ^ n32035 ;
  assign n33675 = n33674 ^ n33389 ;
  assign n33676 = n33391 & ~n33675 ;
  assign n33677 = n33676 ^ n33390 ;
  assign n33345 = n33007 ^ n33006 ;
  assign n33388 = n33387 ^ n33345 ;
  assign n33692 = n33677 ^ n33388 ;
  assign n33693 = ~n32878 & n33692 ;
  assign n33694 = n33693 ^ n33387 ;
  assign n33913 = n33912 ^ n33694 ;
  assign n33914 = n33913 ^ x412 ;
  assign n34123 = n34049 ^ n33914 ;
  assign n34122 = ~n34120 & ~n34121 ;
  assign n34138 = n34123 ^ n34122 ;
  assign n34136 = n33062 & ~n34135 ;
  assign n34137 = n34136 ^ n33059 ;
  assign n34193 = n34138 ^ n34137 ;
  assign n34194 = ~n32815 & ~n34193 ;
  assign n34195 = n34194 ^ n33059 ;
  assign n34190 = n34189 ^ n33062 ;
  assign n34191 = n32390 & ~n34190 ;
  assign n34192 = n34191 ^ n32395 ;
  assign n34262 = n34195 ^ n34192 ;
  assign n34263 = n34262 ^ n34260 ;
  assign n34264 = n34261 & n34263 ;
  assign n34265 = n34264 ^ x102 ;
  assign n34266 = n34265 ^ x101 ;
  assign n34139 = n34138 ^ n34136 ;
  assign n34140 = n34137 & ~n34139 ;
  assign n34141 = n34140 ^ n33059 ;
  assign n34184 = n34141 ^ n33119 ;
  assign n34050 = n34049 ^ n33913 ;
  assign n34051 = ~n33914 & n34050 ;
  assign n34052 = n34051 ^ x412 ;
  assign n33695 = n33694 ^ n32035 ;
  assign n33867 = n33866 ^ n33694 ;
  assign n33868 = n33695 & ~n33867 ;
  assign n33869 = n33868 ^ n32035 ;
  assign n33909 = n33869 ^ n31926 ;
  assign n33344 = n33009 ^ n33008 ;
  assign n33870 = n33462 ^ n33344 ;
  assign n33678 = n33677 ^ n33345 ;
  assign n33679 = n33388 & n33678 ;
  assign n33680 = n33679 ^ n33387 ;
  assign n33871 = n33870 ^ n33680 ;
  assign n33872 = n32972 & ~n33871 ;
  assign n33873 = n33872 ^ n33462 ;
  assign n33910 = n33909 ^ n33873 ;
  assign n33911 = n33910 ^ x411 ;
  assign n34125 = n34052 ^ n33911 ;
  assign n34124 = ~n34122 & ~n34123 ;
  assign n34133 = n34125 ^ n34124 ;
  assign n34185 = n34184 ^ n34133 ;
  assign n34186 = n32808 & ~n34185 ;
  assign n34187 = n34186 ^ n33119 ;
  assign n34267 = n34187 ^ n32403 ;
  assign n34196 = n34195 ^ n34191 ;
  assign n34197 = n34192 & n34196 ;
  assign n34198 = n34197 ^ n32395 ;
  assign n34268 = n34267 ^ n34198 ;
  assign n34269 = n34268 ^ n34265 ;
  assign n34270 = n34266 & n34269 ;
  assign n34271 = n34270 ^ x101 ;
  assign n34272 = n34271 ^ x100 ;
  assign n34199 = n34198 ^ n34187 ;
  assign n34200 = n34198 ^ n32403 ;
  assign n34201 = n34199 & n34200 ;
  assign n34202 = n34201 ^ n32403 ;
  assign n34273 = n34202 ^ n32385 ;
  assign n34053 = n34052 ^ n33910 ;
  assign n34054 = n33911 & ~n34053 ;
  assign n34055 = n34054 ^ x411 ;
  assign n33874 = n33873 ^ n33869 ;
  assign n33681 = n33680 ^ n33344 ;
  assign n33682 = n33011 ^ n33010 ;
  assign n33683 = n33682 ^ n33462 ;
  assign n33684 = n33683 ^ n33344 ;
  assign n33685 = n33684 ^ n33682 ;
  assign n33686 = n33681 & n33685 ;
  assign n33687 = n33686 ^ n33683 ;
  assign n33688 = n33687 ^ n33475 ;
  assign n33689 = n33033 & ~n33688 ;
  assign n33690 = n33689 ^ n33475 ;
  assign n33875 = n33690 ^ n31926 ;
  assign n33876 = n33875 ^ n33869 ;
  assign n33877 = n33876 ^ n33690 ;
  assign n33878 = n33874 & n33877 ;
  assign n33879 = n33878 ^ n33875 ;
  assign n33907 = n33879 ^ n31921 ;
  assign n33908 = n33907 ^ x410 ;
  assign n34127 = n34055 ^ n33908 ;
  assign n34126 = n34124 & n34125 ;
  assign n34145 = n34127 ^ n34126 ;
  assign n34203 = n34145 ^ n33191 ;
  assign n34134 = n34133 ^ n33119 ;
  assign n34142 = n34141 ^ n34133 ;
  assign n34143 = n34134 & ~n34142 ;
  assign n34144 = n34143 ^ n33119 ;
  assign n34204 = n34203 ^ n34144 ;
  assign n34205 = ~n32822 & n34204 ;
  assign n34206 = n34205 ^ n33191 ;
  assign n34274 = n34273 ^ n34206 ;
  assign n34275 = n34274 ^ n34271 ;
  assign n34276 = n34272 & n34275 ;
  assign n34277 = n34276 ^ x100 ;
  assign n34207 = n34206 ^ n34202 ;
  assign n34146 = n34145 ^ n34144 ;
  assign n34128 = ~n34126 & n34127 ;
  assign n33691 = n33690 ^ n31921 ;
  assign n33880 = n33691 & n33879 ;
  assign n33881 = n33880 ^ n31921 ;
  assign n34060 = n33881 ^ n32054 ;
  assign n33884 = n33682 ^ n33475 ;
  assign n33885 = n33687 & ~n33884 ;
  assign n33886 = n33885 ^ n33475 ;
  assign n33882 = n33013 ^ n33012 ;
  assign n33883 = n33882 ^ n33542 ;
  assign n33887 = n33886 ^ n33883 ;
  assign n33888 = n33084 & n33887 ;
  assign n33889 = n33888 ^ n33542 ;
  assign n34061 = n34060 ^ n33889 ;
  assign n34056 = n34055 ^ n33907 ;
  assign n34057 = ~n33908 & n34056 ;
  assign n34058 = n34057 ^ x410 ;
  assign n34059 = n34058 ^ x409 ;
  assign n34065 = n34061 ^ n34059 ;
  assign n34131 = n34128 ^ n34065 ;
  assign n34147 = n34131 ^ n33191 ;
  assign n34148 = n34147 ^ n34131 ;
  assign n34149 = n34148 ^ n34144 ;
  assign n34150 = ~n34146 & ~n34149 ;
  assign n34151 = n34150 ^ n34147 ;
  assign n34180 = n34151 ^ n33772 ;
  assign n34181 = ~n32830 & ~n34180 ;
  assign n34182 = n34181 ^ n33772 ;
  assign n34208 = n34182 ^ n32385 ;
  assign n34209 = n34208 ^ n34182 ;
  assign n34210 = n34209 ^ n34202 ;
  assign n34211 = ~n34207 & ~n34210 ;
  assign n34212 = n34211 ^ n34208 ;
  assign n34257 = n34212 ^ n32382 ;
  assign n34278 = n34277 ^ n34257 ;
  assign n34279 = n34277 ^ x99 ;
  assign n34280 = n34278 & n34279 ;
  assign n34281 = n34280 ^ x99 ;
  assign n34334 = n34281 ^ x98 ;
  assign n34183 = n34182 ^ n32382 ;
  assign n34213 = n34183 & ~n34212 ;
  assign n34214 = n34213 ^ n32382 ;
  assign n34129 = n34065 & n34128 ;
  assign n34062 = n34061 ^ n34058 ;
  assign n34063 = n34059 & n34062 ;
  assign n33900 = n33581 ^ n33014 ;
  assign n33901 = n33900 ^ n33015 ;
  assign n33902 = n33901 ^ n33882 ;
  assign n33897 = n33886 ^ n33882 ;
  assign n33898 = n33886 ^ n33542 ;
  assign n33899 = n33897 & ~n33898 ;
  assign n33903 = n33902 ^ n33899 ;
  assign n33904 = ~n33164 & n33903 ;
  assign n33895 = x409 ^ x408 ;
  assign n33893 = n32069 ^ n32054 ;
  assign n33894 = n33893 ^ n33581 ;
  assign n33896 = n33895 ^ n33894 ;
  assign n33905 = n33904 ^ n33896 ;
  assign n33890 = n33889 ^ n33881 ;
  assign n33891 = n33889 ^ n32054 ;
  assign n33892 = ~n33890 & ~n33891 ;
  assign n33906 = n33905 ^ n33892 ;
  assign n34064 = n34063 ^ n33906 ;
  assign n34130 = n34129 ^ n34064 ;
  assign n34175 = n34130 ^ n33784 ;
  assign n34132 = n34131 ^ n33772 ;
  assign n34152 = ~n34132 & ~n34151 ;
  assign n34153 = n34152 ^ n33772 ;
  assign n34176 = n34175 ^ n34153 ;
  assign n34177 = n32838 & n34176 ;
  assign n34178 = n34177 ^ n33784 ;
  assign n34179 = n34178 ^ n32377 ;
  assign n34255 = n34214 ^ n34179 ;
  assign n34335 = n34334 ^ n34255 ;
  assign n34326 = n34262 ^ n34261 ;
  assign n34327 = n34268 ^ n34266 ;
  assign n34328 = ~n34326 & ~n34327 ;
  assign n34329 = n34274 ^ n34272 ;
  assign n34330 = n34328 & ~n34329 ;
  assign n34331 = n34257 ^ x99 ;
  assign n34332 = n34331 ^ n34277 ;
  assign n34333 = ~n34330 & n34332 ;
  assign n34414 = n34335 ^ n34333 ;
  assign n34356 = n34082 ^ n34081 ;
  assign n34412 = n34356 ^ n33744 ;
  assign n34357 = n34080 ^ n34078 ;
  assign n34358 = n34357 ^ n33823 ;
  assign n34359 = n34077 ^ n34076 ;
  assign n34360 = n34359 ^ n33749 ;
  assign n34364 = n34075 ^ n34074 ;
  assign n34318 = n34073 ^ n34069 ;
  assign n34319 = n34318 ^ n33756 ;
  assign n34243 = n34072 ^ n34070 ;
  assign n34244 = n34243 ^ n33805 ;
  assign n33142 = n33141 ^ n33138 ;
  assign n33337 = n33336 ^ n33142 ;
  assign n33340 = n33140 ^ n33139 ;
  assign n33341 = n33340 ^ n33339 ;
  assign n33343 = n33342 ^ n33139 ;
  assign n34154 = n34153 ^ n34130 ;
  assign n34155 = n33784 ^ n33139 ;
  assign n34156 = n34155 ^ n33139 ;
  assign n34157 = n34156 ^ n34130 ;
  assign n34158 = n34154 & ~n34157 ;
  assign n34159 = n34158 ^ n34155 ;
  assign n34160 = ~n33343 & n34159 ;
  assign n34161 = n34160 ^ n33139 ;
  assign n34162 = n34161 ^ n33339 ;
  assign n34163 = ~n33341 & n34162 ;
  assign n34164 = n34163 ^ n33340 ;
  assign n34165 = n34164 ^ n33336 ;
  assign n34166 = n33337 & n34165 ;
  assign n33202 = n33201 ^ n33200 ;
  assign n33203 = n33202 ^ n33142 ;
  assign n34167 = n34166 ^ n33203 ;
  assign n34240 = n33760 ^ n33202 ;
  assign n34241 = n34167 & ~n34240 ;
  assign n34242 = n34241 ^ n33202 ;
  assign n34315 = n34242 ^ n33805 ;
  assign n34316 = n34244 & n34315 ;
  assign n34317 = n34316 ^ n34243 ;
  assign n34361 = n34317 ^ n33756 ;
  assign n34362 = ~n34319 & ~n34361 ;
  assign n34363 = n34362 ^ n34318 ;
  assign n34365 = n34364 ^ n34363 ;
  assign n34366 = n34359 ^ n33752 ;
  assign n34367 = n34366 ^ n34359 ;
  assign n34368 = n34367 ^ n34363 ;
  assign n34369 = ~n34365 & ~n34368 ;
  assign n34370 = n34369 ^ n34366 ;
  assign n34371 = n34360 & ~n34370 ;
  assign n34372 = n34371 ^ n33749 ;
  assign n34373 = n34372 ^ n34357 ;
  assign n34374 = ~n34358 & ~n34373 ;
  assign n34375 = n34374 ^ n33823 ;
  assign n34413 = n34412 ^ n34375 ;
  assign n34415 = n34414 ^ n34413 ;
  assign n34417 = n34332 ^ n34330 ;
  assign n34854 = n34417 ^ n34413 ;
  assign n34416 = n34372 ^ n34358 ;
  assign n34418 = n34417 ^ n34416 ;
  assign n34420 = n34370 ^ n33749 ;
  assign n34419 = n34329 ^ n34328 ;
  assign n34421 = n34420 ^ n34419 ;
  assign n34843 = n34327 ^ n34326 ;
  assign n34320 = n34319 ^ n34317 ;
  assign n34422 = n34326 ^ n34320 ;
  assign n34423 = n34259 ^ x103 ;
  assign n34245 = n34244 ^ n34242 ;
  assign n34424 = n34423 ^ n34245 ;
  assign n34782 = n33164 ^ n33084 ;
  assign n34783 = n34782 ^ n33903 ;
  assign n34784 = n34783 ^ x120 ;
  assign n34710 = n34116 ^ n34115 ;
  assign n34711 = n34710 ^ n33887 ;
  assign n34461 = n34112 ^ n34111 ;
  assign n34462 = n34461 ^ n33871 ;
  assign n34426 = n34107 ^ n34106 ;
  assign n34427 = n34426 ^ n33696 ;
  assign n34429 = n34098 ^ n34096 ;
  assign n34430 = n34429 ^ n33712 ;
  assign n34399 = n34095 ^ n34067 ;
  assign n34400 = n34399 ^ n33717 ;
  assign n34349 = n34094 ^ n34092 ;
  assign n34350 = n34349 ^ n33722 ;
  assign n34351 = n34091 ^ n34090 ;
  assign n34352 = n34351 ^ n33727 ;
  assign n34353 = n34089 ^ n34087 ;
  assign n34354 = n34353 ^ n33731 ;
  assign n34379 = n33744 ^ n33740 ;
  assign n34376 = n34375 ^ n34356 ;
  assign n34377 = n34375 ^ n33744 ;
  assign n34378 = ~n34376 & ~n34377 ;
  assign n34380 = n34379 ^ n34378 ;
  assign n34381 = n34084 ^ n34083 ;
  assign n34382 = n34381 ^ n33740 ;
  assign n34383 = n34380 & ~n34382 ;
  assign n34355 = n33740 ^ n33735 ;
  assign n34384 = n34383 ^ n34355 ;
  assign n34387 = n34353 ^ n33735 ;
  assign n34385 = n34086 ^ n34085 ;
  assign n34386 = n34385 ^ n34353 ;
  assign n34388 = n34387 ^ n34386 ;
  assign n34389 = n34384 & n34388 ;
  assign n34390 = n34389 ^ n34387 ;
  assign n34391 = n34354 & ~n34390 ;
  assign n34392 = n34391 ^ n33731 ;
  assign n34393 = n34392 ^ n34351 ;
  assign n34394 = ~n34352 & ~n34393 ;
  assign n34395 = n34394 ^ n33727 ;
  assign n34396 = n34395 ^ n34349 ;
  assign n34397 = n34350 & n34396 ;
  assign n34398 = n34397 ^ n33722 ;
  assign n34431 = n34399 ^ n34398 ;
  assign n34432 = n34400 & n34431 ;
  assign n34433 = n34432 ^ n33717 ;
  assign n34434 = n34433 ^ n34429 ;
  assign n34435 = n34430 & n34434 ;
  assign n34436 = n34435 ^ n33712 ;
  assign n34428 = n34100 ^ n34099 ;
  assign n34437 = n34436 ^ n34428 ;
  assign n34438 = n34102 ^ n34101 ;
  assign n34439 = n34438 ^ n33708 ;
  assign n34440 = n34439 ^ n34436 ;
  assign n34441 = n34440 ^ n34438 ;
  assign n34442 = n34437 & ~n34441 ;
  assign n34443 = n34442 ^ n34439 ;
  assign n34444 = n34105 ^ n34103 ;
  assign n34446 = n34444 ^ n33704 ;
  assign n34445 = n34444 ^ n34438 ;
  assign n34447 = n34446 ^ n34445 ;
  assign n34448 = n34443 & n34447 ;
  assign n34449 = n34448 ^ n34446 ;
  assign n34451 = n34426 ^ n33700 ;
  assign n34450 = n34444 ^ n34426 ;
  assign n34452 = n34451 ^ n34450 ;
  assign n34453 = ~n34449 & ~n34452 ;
  assign n34454 = n34453 ^ n34451 ;
  assign n34455 = n34427 & ~n34454 ;
  assign n34456 = n34455 ^ n33696 ;
  assign n34425 = n34110 ^ n34108 ;
  assign n34457 = n34456 ^ n34425 ;
  assign n34458 = n34456 ^ n33692 ;
  assign n34459 = ~n34457 & n34458 ;
  assign n34460 = n34459 ^ n33692 ;
  assign n34589 = n34461 ^ n34460 ;
  assign n34590 = n34462 & n34589 ;
  assign n34591 = n34590 ^ n33871 ;
  assign n34587 = n34114 ^ n34113 ;
  assign n34706 = n34591 ^ n34587 ;
  assign n34707 = n34591 ^ n33688 ;
  assign n34708 = n34706 & n34707 ;
  assign n34709 = n34708 ^ n33688 ;
  assign n34712 = n34711 ^ n34709 ;
  assign n34713 = ~n33542 & ~n34712 ;
  assign n34714 = n34713 ^ n33887 ;
  assign n34715 = n34714 ^ n33084 ;
  assign n34588 = n34587 ^ n33688 ;
  assign n34592 = n34591 ^ n34588 ;
  assign n34593 = ~n33475 & n34592 ;
  assign n34594 = n34593 ^ n33688 ;
  assign n34574 = n34425 ^ n33692 ;
  assign n34575 = n34574 ^ n34456 ;
  assign n34576 = n33387 & n34575 ;
  assign n34577 = n34576 ^ n33692 ;
  assign n34466 = n34454 ^ n33696 ;
  assign n34467 = ~n33390 & n34466 ;
  assign n34468 = n34467 ^ n33696 ;
  assign n34469 = n34468 ^ n32792 ;
  assign n34470 = n34449 ^ n33700 ;
  assign n34471 = ~n33393 & n34470 ;
  assign n34472 = n34471 ^ n33700 ;
  assign n34473 = n34472 ^ n32764 ;
  assign n34560 = n34443 ^ n33704 ;
  assign n34561 = n33397 & n34560 ;
  assign n34562 = n34561 ^ n33704 ;
  assign n34474 = n34437 ^ n33708 ;
  assign n34475 = ~n33399 & ~n34474 ;
  assign n34476 = n34475 ^ n33708 ;
  assign n34477 = n34476 ^ n32327 ;
  assign n34478 = n34433 ^ n34430 ;
  assign n34479 = ~n33411 & n34478 ;
  assign n34480 = n34479 ^ n33712 ;
  assign n34481 = n34480 ^ n32498 ;
  assign n34401 = n34400 ^ n34398 ;
  assign n34482 = ~n33425 & ~n34401 ;
  assign n34483 = n34482 ^ n33717 ;
  assign n34484 = n34483 ^ n32332 ;
  assign n34543 = n34395 ^ n34350 ;
  assign n34544 = ~n33419 & n34543 ;
  assign n34545 = n34544 ^ n33722 ;
  assign n34485 = n34392 ^ n34352 ;
  assign n34486 = n33316 & n34485 ;
  assign n34487 = n34486 ^ n33727 ;
  assign n34488 = n34487 ^ n32336 ;
  assign n34403 = n34390 ^ n33731 ;
  assign n34533 = ~n33297 & ~n34403 ;
  assign n34534 = n34533 ^ n33731 ;
  assign n34406 = n34385 ^ n34384 ;
  assign n34489 = ~n33246 & ~n34406 ;
  assign n34490 = n34489 ^ n33735 ;
  assign n34491 = n34490 ^ n32341 ;
  assign n34409 = n34381 ^ n34380 ;
  assign n34492 = ~n33214 & n34409 ;
  assign n34493 = n34492 ^ n33740 ;
  assign n34494 = n34493 ^ n32465 ;
  assign n34520 = ~n33223 & ~n34413 ;
  assign n34521 = n34520 ^ n33744 ;
  assign n34495 = ~n33175 & n34416 ;
  assign n34496 = n34495 ^ n33823 ;
  assign n34497 = n34496 ^ n32349 ;
  assign n34498 = n33101 & ~n34420 ;
  assign n34499 = n34498 ^ n33749 ;
  assign n34500 = n34499 ^ n32450 ;
  assign n34505 = n34364 ^ n33752 ;
  assign n34506 = n34505 ^ n34363 ;
  assign n34507 = ~n33047 & ~n34506 ;
  assign n34508 = n34507 ^ n33752 ;
  assign n34321 = ~n32985 & n34320 ;
  assign n34322 = n34321 ^ n33756 ;
  assign n34501 = n34322 ^ n32358 ;
  assign n34246 = n32896 & n34245 ;
  assign n34247 = n34246 ^ n33805 ;
  assign n34310 = n34247 ^ n32436 ;
  assign n34168 = n34167 ^ n33760 ;
  assign n34169 = n32801 & ~n34168 ;
  assign n34170 = n34169 ^ n33760 ;
  assign n34171 = n34170 ^ n32362 ;
  assign n34229 = n34164 ^ n33337 ;
  assign n34230 = ~n32861 & ~n34229 ;
  assign n34231 = n34230 ^ n33336 ;
  assign n34222 = n34161 ^ n33341 ;
  assign n34223 = ~n32803 & n34222 ;
  assign n34224 = n34223 ^ n33339 ;
  assign n34215 = n34214 ^ n34178 ;
  assign n34216 = n34179 & ~n34215 ;
  assign n34217 = n34216 ^ n32377 ;
  assign n34172 = n34159 ^ n33342 ;
  assign n34173 = ~n32846 & n34172 ;
  assign n34174 = n34173 ^ n33342 ;
  assign n34218 = n34217 ^ n34174 ;
  assign n34219 = n34217 ^ n32374 ;
  assign n34220 = n34218 & n34219 ;
  assign n34221 = n34220 ^ n32374 ;
  assign n34225 = n34224 ^ n34221 ;
  assign n34226 = n34224 ^ n32369 ;
  assign n34227 = n34225 & n34226 ;
  assign n34228 = n34227 ^ n32369 ;
  assign n34232 = n34231 ^ n34228 ;
  assign n34233 = n34231 ^ n32366 ;
  assign n34234 = ~n34232 & n34233 ;
  assign n34235 = n34234 ^ n32366 ;
  assign n34236 = n34235 ^ n34170 ;
  assign n34237 = ~n34171 & n34236 ;
  assign n34238 = n34237 ^ n32362 ;
  assign n34311 = n34247 ^ n34238 ;
  assign n34312 = ~n34310 & n34311 ;
  assign n34313 = n34312 ^ n32436 ;
  assign n34502 = n34322 ^ n34313 ;
  assign n34503 = ~n34501 & n34502 ;
  assign n34504 = n34503 ^ n32358 ;
  assign n34509 = n34508 ^ n34504 ;
  assign n34510 = n34499 ^ n32353 ;
  assign n34511 = n34510 ^ n34504 ;
  assign n34512 = n34511 ^ n34499 ;
  assign n34513 = n34509 & ~n34512 ;
  assign n34514 = n34513 ^ n34510 ;
  assign n34515 = n34500 & ~n34514 ;
  assign n34516 = n34515 ^ n32450 ;
  assign n34517 = n34516 ^ n34496 ;
  assign n34518 = ~n34497 & n34517 ;
  assign n34519 = n34518 ^ n32349 ;
  assign n34522 = n34521 ^ n34519 ;
  assign n34523 = n34493 ^ n32346 ;
  assign n34524 = n34523 ^ n34493 ;
  assign n34525 = n34524 ^ n34519 ;
  assign n34526 = ~n34522 & ~n34525 ;
  assign n34527 = n34526 ^ n34523 ;
  assign n34528 = ~n34494 & n34527 ;
  assign n34529 = n34528 ^ n32465 ;
  assign n34530 = n34529 ^ n34490 ;
  assign n34531 = ~n34491 & n34530 ;
  assign n34532 = n34531 ^ n32341 ;
  assign n34535 = n34534 ^ n34532 ;
  assign n34536 = n34487 ^ n32475 ;
  assign n34537 = n34536 ^ n34487 ;
  assign n34538 = n34537 ^ n34532 ;
  assign n34539 = n34535 & ~n34538 ;
  assign n34540 = n34539 ^ n34536 ;
  assign n34541 = n34488 & n34540 ;
  assign n34542 = n34541 ^ n32336 ;
  assign n34546 = n34545 ^ n34542 ;
  assign n34547 = n34483 ^ n32486 ;
  assign n34548 = n34547 ^ n34483 ;
  assign n34549 = n34548 ^ n34542 ;
  assign n34550 = n34546 & ~n34549 ;
  assign n34551 = n34550 ^ n34547 ;
  assign n34552 = ~n34484 & n34551 ;
  assign n34553 = n34552 ^ n32332 ;
  assign n34554 = n34553 ^ n34480 ;
  assign n34555 = ~n34481 & ~n34554 ;
  assign n34556 = n34555 ^ n32498 ;
  assign n34557 = n34556 ^ n34476 ;
  assign n34558 = n34477 & ~n34557 ;
  assign n34559 = n34558 ^ n32327 ;
  assign n34563 = n34562 ^ n34559 ;
  assign n34564 = n34472 ^ n32708 ;
  assign n34565 = n34564 ^ n34472 ;
  assign n34566 = n34565 ^ n34559 ;
  assign n34567 = n34563 & ~n34566 ;
  assign n34568 = n34567 ^ n34564 ;
  assign n34569 = ~n34473 & n34568 ;
  assign n34570 = n34569 ^ n32764 ;
  assign n34571 = n34570 ^ n34468 ;
  assign n34572 = ~n34469 & n34571 ;
  assign n34573 = n34572 ^ n32792 ;
  assign n34578 = n34577 ^ n34573 ;
  assign n34579 = n34577 ^ n32878 ;
  assign n34580 = n34578 & ~n34579 ;
  assign n34581 = n34580 ^ n32878 ;
  assign n34463 = n34462 ^ n34460 ;
  assign n34464 = ~n33462 & n34463 ;
  assign n34465 = n34464 ^ n33871 ;
  assign n34582 = n34581 ^ n34465 ;
  assign n34583 = n34581 ^ n32972 ;
  assign n34584 = ~n34582 & ~n34583 ;
  assign n34585 = n34584 ^ n32972 ;
  assign n34702 = n34594 ^ n34585 ;
  assign n34703 = n34594 ^ n33033 ;
  assign n34704 = n34702 & ~n34703 ;
  assign n34705 = n34704 ^ n33033 ;
  assign n34780 = n34714 ^ n34705 ;
  assign n34781 = n34715 & ~n34780 ;
  assign n34785 = n34784 ^ n34781 ;
  assign n34776 = n34709 ^ n33887 ;
  assign n34777 = n34711 & ~n34776 ;
  assign n34773 = n34119 ^ n33903 ;
  assign n34774 = n34773 ^ n34117 ;
  assign n34775 = n34774 ^ n33887 ;
  assign n34778 = n34777 ^ n34775 ;
  assign n34779 = ~n33581 & n34778 ;
  assign n34786 = n34785 ^ n34779 ;
  assign n34695 = n34465 ^ n32972 ;
  assign n34696 = n34695 ^ n34581 ;
  assign n34596 = n34579 ^ n34573 ;
  assign n34597 = n34596 ^ x124 ;
  assign n34598 = n34570 ^ n32792 ;
  assign n34599 = n34598 ^ n34468 ;
  assign n34600 = n34599 ^ x125 ;
  assign n34601 = n34568 ^ n32764 ;
  assign n34602 = n34601 ^ x126 ;
  assign n34603 = n34562 ^ n32708 ;
  assign n34604 = n34603 ^ n34559 ;
  assign n34605 = n34604 ^ x127 ;
  assign n34676 = n34556 ^ n32327 ;
  assign n34677 = n34676 ^ n34476 ;
  assign n34606 = n34553 ^ n32498 ;
  assign n34607 = n34606 ^ n34480 ;
  assign n34608 = n34607 ^ x113 ;
  assign n34609 = n34551 ^ n32332 ;
  assign n34610 = n34609 ^ x114 ;
  assign n34657 = n34540 ^ n32336 ;
  assign n34611 = n34532 ^ n32475 ;
  assign n34612 = n34611 ^ n34534 ;
  assign n34613 = n34612 ^ x117 ;
  assign n34614 = n34529 ^ n34491 ;
  assign n34615 = n34614 ^ x118 ;
  assign n34616 = n34527 ^ n32465 ;
  assign n34617 = n34616 ^ x119 ;
  assign n34641 = n34519 ^ n32346 ;
  assign n34642 = n34641 ^ n34521 ;
  assign n34618 = n34516 ^ n32349 ;
  assign n34619 = n34618 ^ n34496 ;
  assign n34620 = n34619 ^ x105 ;
  assign n34632 = n34514 ^ n32450 ;
  assign n34621 = n34508 ^ n32353 ;
  assign n34622 = n34621 ^ n34504 ;
  assign n34623 = n34622 ^ x107 ;
  assign n34314 = n34313 ^ n32358 ;
  assign n34323 = n34322 ^ n34314 ;
  assign n34239 = n34238 ^ n32436 ;
  assign n34248 = n34247 ^ n34239 ;
  assign n34249 = n34248 ^ x109 ;
  assign n34293 = n34228 ^ n32366 ;
  assign n34294 = n34293 ^ n34231 ;
  assign n34250 = n34221 ^ n32369 ;
  assign n34251 = n34250 ^ n34224 ;
  assign n34252 = n34251 ^ x96 ;
  assign n34256 = n34255 ^ x98 ;
  assign n34282 = n34281 ^ n34255 ;
  assign n34283 = ~n34256 & n34282 ;
  assign n34284 = n34283 ^ x98 ;
  assign n34253 = n34174 ^ n32374 ;
  assign n34254 = n34253 ^ n34217 ;
  assign n34285 = n34284 ^ n34254 ;
  assign n34286 = n34251 ^ x97 ;
  assign n34287 = n34286 ^ n34251 ;
  assign n34288 = n34287 ^ n34254 ;
  assign n34289 = ~n34285 & n34288 ;
  assign n34290 = n34289 ^ n34286 ;
  assign n34291 = ~n34252 & n34290 ;
  assign n34292 = n34291 ^ x96 ;
  assign n34295 = n34294 ^ n34292 ;
  assign n34296 = n34235 ^ n34171 ;
  assign n34297 = n34296 ^ x111 ;
  assign n34298 = n34297 ^ n34292 ;
  assign n34299 = n34298 ^ n34296 ;
  assign n34300 = ~n34295 & n34299 ;
  assign n34301 = n34300 ^ n34297 ;
  assign n34303 = n34248 ^ x110 ;
  assign n34302 = n34296 ^ n34248 ;
  assign n34304 = n34303 ^ n34302 ;
  assign n34305 = n34301 & ~n34304 ;
  assign n34306 = n34305 ^ n34303 ;
  assign n34307 = ~n34249 & n34306 ;
  assign n34308 = n34307 ^ x109 ;
  assign n34624 = n34323 ^ n34308 ;
  assign n34625 = n34622 ^ x108 ;
  assign n34626 = n34625 ^ n34622 ;
  assign n34627 = n34626 ^ n34308 ;
  assign n34628 = n34624 & n34627 ;
  assign n34629 = n34628 ^ n34625 ;
  assign n34630 = n34623 & ~n34629 ;
  assign n34631 = n34630 ^ x107 ;
  assign n34633 = n34632 ^ n34631 ;
  assign n34634 = n34619 ^ x106 ;
  assign n34635 = n34634 ^ n34631 ;
  assign n34636 = n34635 ^ n34619 ;
  assign n34637 = n34633 & n34636 ;
  assign n34638 = n34637 ^ n34634 ;
  assign n34639 = n34620 & ~n34638 ;
  assign n34640 = n34639 ^ x105 ;
  assign n34643 = n34642 ^ n34640 ;
  assign n34644 = n34616 ^ x104 ;
  assign n34645 = n34644 ^ n34616 ;
  assign n34646 = n34645 ^ n34640 ;
  assign n34647 = ~n34643 & n34646 ;
  assign n34648 = n34647 ^ n34644 ;
  assign n34649 = ~n34617 & n34648 ;
  assign n34650 = n34649 ^ x119 ;
  assign n34651 = n34650 ^ n34614 ;
  assign n34652 = ~n34615 & n34651 ;
  assign n34653 = n34652 ^ x118 ;
  assign n34654 = n34653 ^ n34612 ;
  assign n34655 = n34613 & ~n34654 ;
  assign n34656 = n34655 ^ x117 ;
  assign n34658 = n34657 ^ n34656 ;
  assign n34659 = n34545 ^ n32486 ;
  assign n34660 = n34659 ^ n34542 ;
  assign n34661 = n34660 ^ x116 ;
  assign n34662 = n34661 ^ n34656 ;
  assign n34663 = n34662 ^ n34660 ;
  assign n34664 = n34658 & n34663 ;
  assign n34665 = n34664 ^ n34661 ;
  assign n34667 = n34609 ^ x115 ;
  assign n34666 = n34660 ^ n34609 ;
  assign n34668 = n34667 ^ n34666 ;
  assign n34669 = ~n34665 & n34668 ;
  assign n34670 = n34669 ^ n34667 ;
  assign n34671 = n34610 & ~n34670 ;
  assign n34672 = n34671 ^ x114 ;
  assign n34673 = n34672 ^ n34607 ;
  assign n34674 = n34608 & ~n34673 ;
  assign n34675 = n34674 ^ x113 ;
  assign n34678 = n34677 ^ n34675 ;
  assign n34679 = n34604 ^ x112 ;
  assign n34680 = n34679 ^ n34604 ;
  assign n34681 = n34680 ^ n34675 ;
  assign n34682 = ~n34678 & n34681 ;
  assign n34683 = n34682 ^ n34679 ;
  assign n34684 = n34605 & ~n34683 ;
  assign n34685 = n34684 ^ x127 ;
  assign n34686 = n34685 ^ n34601 ;
  assign n34687 = n34602 & ~n34686 ;
  assign n34688 = n34687 ^ x126 ;
  assign n34689 = n34688 ^ n34599 ;
  assign n34690 = n34600 & ~n34689 ;
  assign n34691 = n34690 ^ x125 ;
  assign n34692 = n34691 ^ n34596 ;
  assign n34693 = n34597 & ~n34692 ;
  assign n34694 = n34693 ^ x124 ;
  assign n34697 = n34696 ^ n34694 ;
  assign n34698 = n34696 ^ x123 ;
  assign n34699 = ~n34697 & n34698 ;
  assign n34700 = n34699 ^ x123 ;
  assign n34586 = n34585 ^ n33033 ;
  assign n34595 = n34594 ^ n34586 ;
  assign n34701 = n34700 ^ n34595 ;
  assign n34716 = n34715 ^ n34705 ;
  assign n34717 = n34716 ^ x122 ;
  assign n34718 = n34717 ^ n34595 ;
  assign n34719 = n34718 ^ n34716 ;
  assign n34720 = n34701 & ~n34719 ;
  assign n34721 = n34720 ^ n34717 ;
  assign n34723 = n34700 ^ x122 ;
  assign n34724 = n34723 ^ n34595 ;
  assign n34725 = n34698 ^ n34694 ;
  assign n34726 = n34632 ^ x106 ;
  assign n34727 = n34726 ^ n34631 ;
  assign n34309 = n34308 ^ x108 ;
  assign n34324 = n34323 ^ n34309 ;
  assign n34325 = n34301 ^ x110 ;
  assign n34336 = ~n34333 & ~n34335 ;
  assign n34337 = n34254 ^ x97 ;
  assign n34338 = n34337 ^ n34284 ;
  assign n34339 = n34336 & n34338 ;
  assign n34340 = n34290 ^ x96 ;
  assign n34341 = ~n34339 & n34340 ;
  assign n34342 = n34294 ^ x111 ;
  assign n34343 = n34342 ^ n34292 ;
  assign n34344 = ~n34341 & n34343 ;
  assign n34345 = ~n34325 & n34344 ;
  assign n34346 = n34306 ^ x109 ;
  assign n34347 = ~n34345 & n34346 ;
  assign n34728 = n34324 & n34347 ;
  assign n34729 = n34629 ^ x107 ;
  assign n34730 = ~n34728 & n34729 ;
  assign n34731 = ~n34727 & n34730 ;
  assign n34732 = n34638 ^ x105 ;
  assign n34733 = ~n34731 & ~n34732 ;
  assign n34734 = n34642 ^ x104 ;
  assign n34735 = n34734 ^ n34640 ;
  assign n34736 = n34733 & ~n34735 ;
  assign n34737 = n34648 ^ x119 ;
  assign n34738 = ~n34736 & ~n34737 ;
  assign n34739 = n34650 ^ x118 ;
  assign n34740 = n34739 ^ n34614 ;
  assign n34741 = n34738 & ~n34740 ;
  assign n34742 = n34653 ^ n34613 ;
  assign n34743 = ~n34741 & ~n34742 ;
  assign n34744 = n34657 ^ x116 ;
  assign n34745 = n34744 ^ n34656 ;
  assign n34746 = n34743 & n34745 ;
  assign n34747 = n34665 ^ x115 ;
  assign n34748 = ~n34746 & n34747 ;
  assign n34749 = n34670 ^ x114 ;
  assign n34750 = n34748 & n34749 ;
  assign n34751 = n34672 ^ x113 ;
  assign n34752 = n34751 ^ n34607 ;
  assign n34753 = n34750 & n34752 ;
  assign n34754 = n34677 ^ x112 ;
  assign n34755 = n34754 ^ n34675 ;
  assign n34756 = n34753 & n34755 ;
  assign n34757 = n34683 ^ x127 ;
  assign n34758 = ~n34756 & ~n34757 ;
  assign n34759 = n34685 ^ x126 ;
  assign n34760 = n34759 ^ n34601 ;
  assign n34761 = n34758 & ~n34760 ;
  assign n34762 = n34688 ^ n34600 ;
  assign n34763 = n34761 & ~n34762 ;
  assign n34764 = n34691 ^ n34597 ;
  assign n34765 = n34763 & ~n34764 ;
  assign n34766 = n34725 & ~n34765 ;
  assign n34767 = ~n34724 & n34766 ;
  assign n34768 = n34767 ^ n34716 ;
  assign n34771 = ~n34721 & ~n34768 ;
  assign n34722 = n34721 ^ n34716 ;
  assign n34769 = n34768 ^ n34722 ;
  assign n34770 = ~x121 & n34769 ;
  assign n34772 = n34771 ^ n34770 ;
  assign n34787 = n34786 ^ n34772 ;
  assign n34788 = n34787 ^ n34168 ;
  assign n34821 = n34766 ^ n34724 ;
  assign n34789 = n34765 ^ n34725 ;
  assign n34790 = n34789 ^ n34172 ;
  assign n34791 = n34764 ^ n34763 ;
  assign n34792 = n34791 ^ n34176 ;
  assign n34793 = n34762 ^ n34761 ;
  assign n34794 = n34793 ^ n34180 ;
  assign n34795 = n34760 ^ n34758 ;
  assign n34796 = n34795 ^ n34204 ;
  assign n34797 = n34752 ^ n34750 ;
  assign n34798 = ~n34188 & n34797 ;
  assign n34799 = n34798 ^ n34193 ;
  assign n34800 = n34755 ^ n34753 ;
  assign n34801 = n34800 ^ n34798 ;
  assign n34802 = n34799 & ~n34801 ;
  assign n34803 = n34802 ^ n34193 ;
  assign n34804 = n34803 ^ n34185 ;
  assign n34805 = n34757 ^ n34756 ;
  assign n34806 = n34805 ^ n34803 ;
  assign n34807 = n34804 & n34806 ;
  assign n34808 = n34807 ^ n34185 ;
  assign n34809 = n34808 ^ n34795 ;
  assign n34810 = ~n34796 & ~n34809 ;
  assign n34811 = n34810 ^ n34204 ;
  assign n34812 = n34811 ^ n34793 ;
  assign n34813 = n34794 & n34812 ;
  assign n34814 = n34813 ^ n34180 ;
  assign n34815 = n34814 ^ n34791 ;
  assign n34816 = ~n34792 & ~n34815 ;
  assign n34817 = n34816 ^ n34176 ;
  assign n34818 = n34817 ^ n34789 ;
  assign n34819 = n34790 & ~n34818 ;
  assign n34820 = n34819 ^ n34172 ;
  assign n34822 = n34821 ^ n34820 ;
  assign n34823 = n34721 ^ x121 ;
  assign n34824 = n34823 ^ n34767 ;
  assign n34825 = n34824 ^ n34222 ;
  assign n34826 = n34825 ^ n34820 ;
  assign n34827 = n34826 ^ n34824 ;
  assign n34828 = ~n34822 & n34827 ;
  assign n34829 = n34828 ^ n34825 ;
  assign n34831 = n34787 ^ n34229 ;
  assign n34830 = n34824 ^ n34787 ;
  assign n34832 = n34831 ^ n34830 ;
  assign n34833 = n34829 & n34832 ;
  assign n34834 = n34833 ^ n34831 ;
  assign n34835 = ~n34788 & n34834 ;
  assign n34836 = n34835 ^ n34168 ;
  assign n34837 = n34836 ^ n34423 ;
  assign n34838 = n34424 & n34837 ;
  assign n34839 = n34838 ^ n34245 ;
  assign n34840 = n34839 ^ n34326 ;
  assign n34841 = ~n34422 & n34840 ;
  assign n34842 = n34841 ^ n34320 ;
  assign n34844 = n34843 ^ n34842 ;
  assign n34847 = n34842 ^ n34506 ;
  assign n34848 = n34844 & ~n34847 ;
  assign n34845 = n34506 ^ n34420 ;
  assign n34849 = n34848 ^ n34845 ;
  assign n34850 = ~n34421 & n34849 ;
  assign n34851 = n34850 ^ n34420 ;
  assign n34852 = n34851 ^ n34416 ;
  assign n34853 = ~n34418 & n34852 ;
  assign n34855 = n34854 ^ n34853 ;
  assign n34856 = n34415 & ~n34855 ;
  assign n34857 = n34856 ^ n34414 ;
  assign n34410 = n34338 ^ n34336 ;
  assign n34411 = n34410 ^ n34409 ;
  assign n35107 = n34857 ^ n34411 ;
  assign n35108 = n33740 & n35107 ;
  assign n35109 = n35108 ^ n34409 ;
  assign n35111 = n35109 ^ n33214 ;
  assign n35038 = n34855 ^ n34414 ;
  assign n35039 = n33744 & ~n35038 ;
  assign n35040 = n35039 ^ n34413 ;
  assign n35041 = n35040 ^ n33223 ;
  assign n35097 = n34851 ^ n34418 ;
  assign n35098 = ~n33823 & n35097 ;
  assign n35099 = n35098 ^ n34416 ;
  assign n35042 = n34843 ^ n34506 ;
  assign n35043 = n35042 ^ n34842 ;
  assign n35044 = n33752 & n35043 ;
  assign n35045 = n35044 ^ n34506 ;
  assign n35046 = n35045 ^ n33047 ;
  assign n35080 = n34839 ^ n34422 ;
  assign n35081 = n33756 & ~n35080 ;
  assign n35082 = n35081 ^ n34320 ;
  assign n35047 = n34836 ^ n34424 ;
  assign n35048 = n33805 & ~n35047 ;
  assign n35049 = n35048 ^ n34245 ;
  assign n35050 = n35049 ^ n32896 ;
  assign n35065 = n34829 ^ n34229 ;
  assign n35066 = ~n33336 & n35065 ;
  assign n35067 = n35066 ^ n34229 ;
  assign n35054 = n34820 ^ n34222 ;
  assign n35055 = n35054 ^ n34821 ;
  assign n35056 = ~n33339 & n35055 ;
  assign n35057 = n35056 ^ n34222 ;
  assign n35058 = n35057 ^ n32803 ;
  assign n34888 = n34814 ^ n34792 ;
  assign n34889 = n33784 & n34888 ;
  assign n34890 = n34889 ^ n34176 ;
  assign n34891 = n34890 ^ n32838 ;
  assign n34892 = n34811 ^ n34794 ;
  assign n34893 = n33772 & n34892 ;
  assign n34894 = n34893 ^ n34180 ;
  assign n34895 = n34894 ^ n32830 ;
  assign n34896 = n34808 ^ n34796 ;
  assign n34897 = ~n33191 & n34896 ;
  assign n34898 = n34897 ^ n34204 ;
  assign n34899 = n34898 ^ n32822 ;
  assign n34903 = n34797 ^ n34135 ;
  assign n34904 = n34903 ^ n33062 ;
  assign n34905 = n33062 & n34904 ;
  assign n34906 = n34905 ^ n34188 ;
  assign n34907 = n32802 & n34906 ;
  assign n34908 = n34907 ^ n32815 ;
  assign n34909 = n34800 ^ n34799 ;
  assign n34910 = n33059 & ~n34909 ;
  assign n34911 = n34910 ^ n34193 ;
  assign n34912 = n34911 ^ n34907 ;
  assign n34913 = ~n34908 & n34912 ;
  assign n34914 = n34913 ^ n32815 ;
  assign n34900 = n34805 ^ n34804 ;
  assign n34901 = n33119 & n34900 ;
  assign n34902 = n34901 ^ n34185 ;
  assign n34915 = n34914 ^ n34902 ;
  assign n34916 = n34914 ^ n32808 ;
  assign n34917 = ~n34915 & ~n34916 ;
  assign n34918 = n34917 ^ n32808 ;
  assign n34919 = n34918 ^ n34898 ;
  assign n34920 = ~n34899 & ~n34919 ;
  assign n34921 = n34920 ^ n32822 ;
  assign n34922 = n34921 ^ n34894 ;
  assign n34923 = n34895 & ~n34922 ;
  assign n34924 = n34923 ^ n32830 ;
  assign n34925 = n34924 ^ n34890 ;
  assign n34926 = n34891 & n34925 ;
  assign n34927 = n34926 ^ n32838 ;
  assign n34928 = n34927 ^ n32846 ;
  assign n34885 = n34817 ^ n34790 ;
  assign n34886 = ~n33342 & n34885 ;
  assign n34887 = n34886 ^ n34172 ;
  assign n35059 = n34927 ^ n34887 ;
  assign n35060 = ~n34928 & ~n35059 ;
  assign n35061 = n35060 ^ n32846 ;
  assign n35062 = n35061 ^ n35057 ;
  assign n35063 = ~n35058 & n35062 ;
  assign n35064 = n35063 ^ n32803 ;
  assign n35068 = n35067 ^ n35064 ;
  assign n35069 = n35067 ^ n32861 ;
  assign n35070 = ~n35068 & n35069 ;
  assign n35071 = n35070 ^ n32861 ;
  assign n35051 = n34834 ^ n34168 ;
  assign n35052 = n33760 & n35051 ;
  assign n35053 = n35052 ^ n34168 ;
  assign n35072 = n35071 ^ n35053 ;
  assign n35073 = n35049 ^ n32801 ;
  assign n35074 = n35073 ^ n35049 ;
  assign n35075 = n35074 ^ n35053 ;
  assign n35076 = ~n35072 & ~n35075 ;
  assign n35077 = n35076 ^ n35073 ;
  assign n35078 = n35050 & ~n35077 ;
  assign n35079 = n35078 ^ n32896 ;
  assign n35083 = n35082 ^ n35079 ;
  assign n35084 = n35082 ^ n32985 ;
  assign n35085 = ~n35083 & ~n35084 ;
  assign n35086 = n35085 ^ n32985 ;
  assign n35087 = n35086 ^ n35045 ;
  assign n35088 = n35046 & ~n35087 ;
  assign n35089 = n35088 ^ n33047 ;
  assign n35090 = n35089 ^ n33101 ;
  assign n35091 = n34849 ^ n34419 ;
  assign n35092 = n33749 & n35091 ;
  assign n35093 = n35092 ^ n34420 ;
  assign n35094 = n35093 ^ n35089 ;
  assign n35095 = ~n35090 & ~n35094 ;
  assign n35096 = n35095 ^ n33101 ;
  assign n35100 = n35099 ^ n35096 ;
  assign n35101 = n35099 ^ n33175 ;
  assign n35102 = ~n35100 & ~n35101 ;
  assign n35103 = n35102 ^ n33175 ;
  assign n35104 = n35103 ^ n35040 ;
  assign n35105 = n35041 & ~n35104 ;
  assign n35106 = n35105 ^ n33223 ;
  assign n35266 = n35111 ^ n35106 ;
  assign n35216 = n35103 ^ n35041 ;
  assign n35217 = n35216 ^ x328 ;
  assign n35218 = n35093 ^ n35090 ;
  assign n35219 = n35218 ^ x330 ;
  assign n35220 = n35086 ^ n35046 ;
  assign n35221 = n35220 ^ x331 ;
  assign n35246 = n35084 ^ n35079 ;
  assign n35222 = n35071 ^ n32801 ;
  assign n35223 = n35222 ^ n35053 ;
  assign n35224 = n35223 ^ x334 ;
  assign n34930 = n34924 ^ n34891 ;
  assign n34931 = n34930 ^ x322 ;
  assign n34932 = n34921 ^ n34895 ;
  assign n34933 = n34932 ^ x323 ;
  assign n34936 = n34135 ^ n33017 ;
  assign n34937 = n34936 ^ n34905 ;
  assign n34938 = x327 & n34937 ;
  assign n34939 = n34938 ^ x326 ;
  assign n34940 = n34911 ^ n34908 ;
  assign n34941 = n34940 ^ n34938 ;
  assign n34942 = n34939 & ~n34941 ;
  assign n34943 = n34942 ^ x326 ;
  assign n34944 = n34943 ^ x325 ;
  assign n34945 = n34902 ^ n32808 ;
  assign n34946 = n34945 ^ n34914 ;
  assign n34947 = n34946 ^ n34943 ;
  assign n34948 = n34944 & ~n34947 ;
  assign n34949 = n34948 ^ x325 ;
  assign n34934 = n34918 ^ n32822 ;
  assign n34935 = n34934 ^ n34898 ;
  assign n34950 = n34949 ^ n34935 ;
  assign n34951 = n34949 ^ x324 ;
  assign n34952 = n34950 & n34951 ;
  assign n34953 = n34952 ^ x324 ;
  assign n34954 = n34953 ^ n34932 ;
  assign n34955 = ~n34933 & n34954 ;
  assign n34956 = n34955 ^ x323 ;
  assign n34957 = n34956 ^ n34930 ;
  assign n34958 = ~n34931 & n34957 ;
  assign n34959 = n34958 ^ x322 ;
  assign n34960 = n34959 ^ x321 ;
  assign n34929 = n34928 ^ n34887 ;
  assign n35225 = n34959 ^ n34929 ;
  assign n35226 = n34960 & n35225 ;
  assign n35227 = n35226 ^ x321 ;
  assign n35228 = n35227 ^ x320 ;
  assign n35229 = n35061 ^ n35058 ;
  assign n35230 = n35229 ^ n35227 ;
  assign n35231 = n35228 & ~n35230 ;
  assign n35232 = n35231 ^ x320 ;
  assign n35233 = n35232 ^ x335 ;
  assign n35234 = n35069 ^ n35064 ;
  assign n35235 = n35234 ^ n35232 ;
  assign n35236 = n35233 & n35235 ;
  assign n35237 = n35236 ^ x335 ;
  assign n35238 = n35237 ^ n35223 ;
  assign n35239 = n35224 & ~n35238 ;
  assign n35240 = n35239 ^ x334 ;
  assign n35241 = n35240 ^ x333 ;
  assign n35242 = n35077 ^ n32896 ;
  assign n35243 = n35242 ^ n35240 ;
  assign n35244 = n35241 & ~n35243 ;
  assign n35245 = n35244 ^ x333 ;
  assign n35247 = n35246 ^ n35245 ;
  assign n35248 = n35220 ^ x332 ;
  assign n35249 = n35248 ^ n35220 ;
  assign n35250 = n35249 ^ n35245 ;
  assign n35251 = n35247 & n35250 ;
  assign n35252 = n35251 ^ n35248 ;
  assign n35253 = ~n35221 & n35252 ;
  assign n35254 = n35253 ^ x331 ;
  assign n35255 = n35254 ^ n35218 ;
  assign n35256 = n35219 & ~n35255 ;
  assign n35257 = n35256 ^ x330 ;
  assign n35258 = n35257 ^ x329 ;
  assign n35259 = n35101 ^ n35096 ;
  assign n35260 = n35259 ^ n35257 ;
  assign n35261 = n35258 & n35260 ;
  assign n35262 = n35261 ^ x329 ;
  assign n35263 = n35262 ^ n35216 ;
  assign n35264 = ~n35217 & n35263 ;
  assign n35265 = n35264 ^ x328 ;
  assign n35267 = n35266 ^ n35265 ;
  assign n35268 = n35266 ^ x343 ;
  assign n35269 = ~n35267 & n35268 ;
  assign n35270 = n35269 ^ x343 ;
  assign n35110 = n35109 ^ n35106 ;
  assign n35112 = n35110 & ~n35111 ;
  assign n35113 = n35112 ^ n33214 ;
  assign n35213 = n35113 ^ n33246 ;
  assign n34860 = n34410 ^ n34406 ;
  assign n34858 = n34857 ^ n34409 ;
  assign n34859 = ~n34411 & n34858 ;
  assign n34861 = n34860 ^ n34859 ;
  assign n34407 = n34340 ^ n34339 ;
  assign n34985 = n34861 ^ n34407 ;
  assign n35035 = n33735 & ~n34985 ;
  assign n35036 = n35035 ^ n34406 ;
  assign n35214 = n35213 ^ n35036 ;
  assign n35215 = n35214 ^ x342 ;
  assign n35344 = n35270 ^ n35215 ;
  assign n34961 = n34960 ^ n34929 ;
  assign n34962 = n34956 ^ n34931 ;
  assign n34963 = n34937 ^ x327 ;
  assign n34964 = n34940 ^ n34939 ;
  assign n34965 = n34963 & n34964 ;
  assign n34966 = n34946 ^ n34944 ;
  assign n34967 = ~n34965 & ~n34966 ;
  assign n34968 = n34935 ^ x324 ;
  assign n34969 = n34968 ^ n34949 ;
  assign n34970 = n34967 & n34969 ;
  assign n34971 = n34953 ^ n34933 ;
  assign n34972 = n34970 & n34971 ;
  assign n34973 = n34962 & n34972 ;
  assign n35322 = n34961 & n34973 ;
  assign n35323 = n35229 ^ n35228 ;
  assign n35324 = ~n35322 & n35323 ;
  assign n35325 = n35234 ^ n35233 ;
  assign n35326 = n35324 & ~n35325 ;
  assign n35327 = n35237 ^ n35224 ;
  assign n35328 = n35326 & n35327 ;
  assign n35329 = n35242 ^ n35241 ;
  assign n35330 = ~n35328 & ~n35329 ;
  assign n35331 = n35246 ^ x332 ;
  assign n35332 = n35331 ^ n35245 ;
  assign n35333 = ~n35330 & ~n35332 ;
  assign n35334 = n35252 ^ x331 ;
  assign n35335 = ~n35333 & n35334 ;
  assign n35336 = n35254 ^ n35219 ;
  assign n35337 = n35335 & ~n35336 ;
  assign n35338 = n35259 ^ n35258 ;
  assign n35339 = n35337 & n35338 ;
  assign n35340 = n35262 ^ n35217 ;
  assign n35341 = n35339 & n35340 ;
  assign n35342 = n35268 ^ n35265 ;
  assign n35343 = n35341 & ~n35342 ;
  assign n35395 = n35344 ^ n35343 ;
  assign n35509 = n35395 ^ n34904 ;
  assign n35510 = ~n34188 & ~n35509 ;
  assign n35511 = n35510 ^ n34903 ;
  assign n35512 = n35511 ^ x39 ;
  assign n35271 = n35270 ^ n35214 ;
  assign n35272 = ~n35215 & n35271 ;
  assign n35273 = n35272 ^ x342 ;
  assign n34408 = n34407 ^ n34406 ;
  assign n34862 = n34408 & ~n34861 ;
  assign n34863 = n34862 ^ n34407 ;
  assign n34404 = n34343 ^ n34341 ;
  assign n34405 = n34404 ^ n34403 ;
  assign n34982 = n34863 ^ n34405 ;
  assign n35118 = n33731 & n34982 ;
  assign n35119 = n35118 ^ n34403 ;
  assign n35037 = n35036 ^ n33246 ;
  assign n35114 = n35113 ^ n35036 ;
  assign n35115 = n35037 & ~n35114 ;
  assign n35116 = n35115 ^ n33246 ;
  assign n35117 = n35116 ^ n33297 ;
  assign n35211 = n35119 ^ n35117 ;
  assign n35212 = n35211 ^ x341 ;
  assign n35346 = n35273 ^ n35212 ;
  assign n35345 = n35343 & n35344 ;
  assign n35398 = n35346 ^ n35345 ;
  assign n35396 = ~n34904 & ~n35395 ;
  assign n35399 = n35398 ^ n35396 ;
  assign n35591 = n35399 ^ n34909 ;
  assign n35592 = n34193 & n35591 ;
  assign n35593 = n35592 ^ n34909 ;
  assign n35589 = n33062 & ~n35511 ;
  assign n35590 = n35589 ^ n33059 ;
  assign n35722 = n35593 ^ n35590 ;
  assign n35720 = x39 & n35511 ;
  assign n35721 = n35720 ^ x38 ;
  assign n35852 = n35722 ^ n35721 ;
  assign n35853 = n35512 & ~n35852 ;
  assign n35397 = n35396 ^ n34909 ;
  assign n35400 = n35397 & n35399 ;
  assign n35401 = n35400 ^ n34909 ;
  assign n35599 = n35401 ^ n34900 ;
  assign n35274 = n35273 ^ n35211 ;
  assign n35275 = ~n35212 & n35274 ;
  assign n35276 = n35275 ^ x341 ;
  assign n34870 = n34344 ^ n34325 ;
  assign n34866 = n34485 ^ n34404 ;
  assign n34864 = n34863 ^ n34403 ;
  assign n34865 = ~n34405 & ~n34864 ;
  assign n34867 = n34866 ^ n34865 ;
  assign n35124 = n34870 ^ n34867 ;
  assign n35125 = ~n33727 & n35124 ;
  assign n35126 = n35125 ^ n34485 ;
  assign n35120 = n35119 ^ n35116 ;
  assign n35121 = n35117 & ~n35120 ;
  assign n35122 = n35121 ^ n33297 ;
  assign n35123 = n35122 ^ n33316 ;
  assign n35209 = n35126 ^ n35123 ;
  assign n35210 = n35209 ^ x340 ;
  assign n35348 = n35276 ^ n35210 ;
  assign n35347 = n35345 & n35346 ;
  assign n35402 = n35348 ^ n35347 ;
  assign n35600 = n35599 ^ n35402 ;
  assign n35601 = n34185 & ~n35600 ;
  assign n35594 = n35593 ^ n35589 ;
  assign n35595 = n35590 & n35594 ;
  assign n35596 = n35595 ^ n33059 ;
  assign n35598 = n35596 ^ n34900 ;
  assign n35602 = n35601 ^ n35598 ;
  assign n35727 = n35602 ^ n33119 ;
  assign n35723 = n35722 ^ n35720 ;
  assign n35724 = n35721 & n35723 ;
  assign n35725 = n35724 ^ x38 ;
  assign n35726 = n35725 ^ x37 ;
  assign n35854 = n35727 ^ n35726 ;
  assign n35855 = n35853 & n35854 ;
  assign n35728 = n35727 ^ n35725 ;
  assign n35729 = n35726 & ~n35728 ;
  assign n35730 = n35729 ^ x37 ;
  assign n35856 = n35730 ^ x36 ;
  assign n35597 = n35596 ^ n33119 ;
  assign n35603 = n35597 & ~n35602 ;
  assign n35604 = n35603 ^ n33119 ;
  assign n35403 = n35402 ^ n35401 ;
  assign n35277 = n35276 ^ n35209 ;
  assign n35278 = ~n35210 & n35277 ;
  assign n35279 = n35278 ^ x340 ;
  assign n34868 = n34346 ^ n34345 ;
  assign n34871 = n34870 ^ n34868 ;
  assign n34869 = n34868 ^ n34485 ;
  assign n34872 = n34871 ^ n34869 ;
  assign n34873 = ~n34867 & n34872 ;
  assign n34874 = n34873 ^ n34871 ;
  assign n34978 = n34874 ^ n34543 ;
  assign n35033 = n33722 & ~n34978 ;
  assign n35034 = n35033 ^ n34543 ;
  assign n35206 = n35034 ^ n33419 ;
  assign n35127 = n35126 ^ n35122 ;
  assign n35128 = ~n35123 & n35127 ;
  assign n35129 = n35128 ^ n33316 ;
  assign n35207 = n35206 ^ n35129 ;
  assign n35208 = n35207 ^ x339 ;
  assign n35350 = n35279 ^ n35208 ;
  assign n35349 = n35347 & n35348 ;
  assign n35393 = n35350 ^ n35349 ;
  assign n35404 = n35393 ^ n34900 ;
  assign n35405 = n35404 ^ n35393 ;
  assign n35406 = n35405 ^ n35401 ;
  assign n35407 = n35403 & ~n35406 ;
  assign n35408 = n35407 ^ n35404 ;
  assign n35585 = n35408 ^ n34896 ;
  assign n35586 = ~n34204 & ~n35585 ;
  assign n35587 = n35586 ^ n34896 ;
  assign n35588 = n35587 ^ n33191 ;
  assign n35731 = n35604 ^ n35588 ;
  assign n35857 = n35856 ^ n35731 ;
  assign n35858 = n35855 & ~n35857 ;
  assign n35732 = n35731 ^ n35730 ;
  assign n35736 = n35732 & n35856 ;
  assign n35130 = n35129 ^ n35034 ;
  assign n34348 = n34347 ^ n34324 ;
  assign n34876 = n34543 ^ n34348 ;
  assign n34875 = n34868 ^ n34348 ;
  assign n34877 = n34876 ^ n34875 ;
  assign n34878 = n34874 & ~n34877 ;
  assign n34879 = n34878 ^ n34876 ;
  assign n34975 = n34879 ^ n34401 ;
  assign n35030 = ~n33717 & ~n34975 ;
  assign n35031 = n35030 ^ n34401 ;
  assign n35131 = n35031 ^ n33419 ;
  assign n35132 = n35131 ^ n35031 ;
  assign n35133 = n35132 ^ n35034 ;
  assign n35134 = ~n35130 & ~n35133 ;
  assign n35135 = n35134 ^ n35131 ;
  assign n35284 = n35135 ^ n33425 ;
  assign n35280 = n35279 ^ n35207 ;
  assign n35281 = ~n35208 & n35280 ;
  assign n35282 = n35281 ^ x339 ;
  assign n35283 = n35282 ^ x338 ;
  assign n35352 = n35284 ^ n35283 ;
  assign n35351 = ~n35349 & ~n35350 ;
  assign n35412 = n35352 ^ n35351 ;
  assign n35394 = n35393 ^ n34896 ;
  assign n35409 = ~n35394 & n35408 ;
  assign n35410 = n35409 ^ n34896 ;
  assign n35411 = n35410 ^ n34892 ;
  assign n35609 = n35412 ^ n35411 ;
  assign n35610 = n34180 & ~n35609 ;
  assign n35605 = n35604 ^ n35587 ;
  assign n35606 = ~n35588 & ~n35605 ;
  assign n35607 = n35606 ^ n33191 ;
  assign n35608 = n35607 ^ n34892 ;
  assign n35611 = n35610 ^ n35608 ;
  assign n35718 = n35611 ^ n33772 ;
  assign n35733 = n35718 ^ x36 ;
  assign n35737 = n35736 ^ n35733 ;
  assign n35859 = n35737 ^ x35 ;
  assign n35860 = ~n35858 & n35859 ;
  assign n35413 = n35412 ^ n35410 ;
  assign n35414 = n35411 & n35413 ;
  assign n35415 = n35414 ^ n34892 ;
  assign n35580 = n35415 ^ n34888 ;
  assign n35285 = n35284 ^ n35282 ;
  assign n35286 = n35283 & n35285 ;
  assign n35287 = n35286 ^ x338 ;
  assign n35354 = n35287 ^ x337 ;
  assign n34882 = n34729 ^ n34728 ;
  assign n34883 = n34882 ^ n34478 ;
  assign n34402 = n34401 ^ n34348 ;
  assign n34880 = ~n34402 & ~n34879 ;
  assign n34881 = n34880 ^ n34401 ;
  assign n34884 = n34883 ^ n34881 ;
  assign n35138 = n33712 & ~n34884 ;
  assign n35139 = n35138 ^ n34478 ;
  assign n35141 = n35139 ^ n33411 ;
  assign n35032 = n35031 ^ n33425 ;
  assign n35136 = n35032 & ~n35135 ;
  assign n35137 = n35136 ^ n33425 ;
  assign n35288 = n35141 ^ n35137 ;
  assign n35355 = n35354 ^ n35288 ;
  assign n35353 = ~n35351 & n35352 ;
  assign n35391 = n35355 ^ n35353 ;
  assign n35581 = n35580 ^ n35391 ;
  assign n35582 = ~n34176 & ~n35581 ;
  assign n35583 = n35582 ^ n34888 ;
  assign n35613 = n35583 ^ n33772 ;
  assign n35612 = n35607 ^ n35583 ;
  assign n35614 = n35613 ^ n35612 ;
  assign n35615 = n35611 & ~n35614 ;
  assign n35616 = n35615 ^ n35613 ;
  assign n35741 = n35616 ^ n33784 ;
  assign n35719 = n35718 ^ x35 ;
  assign n35738 = ~n35719 & n35737 ;
  assign n35739 = n35738 ^ x35 ;
  assign n35740 = n35739 ^ x34 ;
  assign n35861 = n35741 ^ n35740 ;
  assign n35862 = ~n35860 & n35861 ;
  assign n35742 = n35741 ^ n35739 ;
  assign n35743 = n35740 & ~n35742 ;
  assign n35744 = n35743 ^ x34 ;
  assign n35584 = n35583 ^ n33784 ;
  assign n35617 = n35584 & ~n35616 ;
  assign n35618 = n35617 ^ n33784 ;
  assign n35392 = n35391 ^ n34888 ;
  assign n35416 = n35415 ^ n35391 ;
  assign n35417 = ~n35392 & n35416 ;
  assign n35418 = n35417 ^ n34888 ;
  assign n35575 = n35418 ^ n34885 ;
  assign n35289 = n35288 ^ n35287 ;
  assign n35140 = n35139 ^ n35137 ;
  assign n35142 = n35140 & ~n35141 ;
  assign n35143 = n35142 ^ n33411 ;
  assign n35203 = n35143 ^ n33399 ;
  assign n34992 = n34881 ^ n34478 ;
  assign n34993 = n34883 & n34992 ;
  assign n34994 = n34993 ^ n34882 ;
  assign n34990 = n34730 ^ n34727 ;
  assign n34991 = n34990 ^ n34474 ;
  assign n35026 = n34994 ^ n34991 ;
  assign n35027 = ~n33708 & ~n35026 ;
  assign n35028 = n35027 ^ n34474 ;
  assign n35204 = n35203 ^ n35028 ;
  assign n35290 = n35204 ^ x337 ;
  assign n35291 = n35290 ^ n35204 ;
  assign n35292 = n35291 ^ n35287 ;
  assign n35293 = ~n35289 & n35292 ;
  assign n35294 = n35293 ^ n35290 ;
  assign n35357 = n35294 ^ x336 ;
  assign n35356 = n35353 & ~n35355 ;
  assign n35389 = n35357 ^ n35356 ;
  assign n35576 = n35575 ^ n35389 ;
  assign n35577 = ~n34172 & n35576 ;
  assign n35578 = n35577 ^ n34885 ;
  assign n35579 = n35578 ^ n33342 ;
  assign n35716 = n35618 ^ n35579 ;
  assign n35717 = n35716 ^ x33 ;
  assign n35863 = n35744 ^ n35717 ;
  assign n35864 = ~n35862 & n35863 ;
  assign n35745 = n35744 ^ n35716 ;
  assign n35746 = ~n35717 & n35745 ;
  assign n35747 = n35746 ^ x33 ;
  assign n35619 = n35618 ^ n35578 ;
  assign n35620 = ~n35579 & ~n35619 ;
  assign n35621 = n35620 ^ n33342 ;
  assign n35358 = n35356 & n35357 ;
  assign n35205 = n35204 ^ x336 ;
  assign n35295 = ~n35205 & n35294 ;
  assign n35296 = n35295 ^ x336 ;
  assign n34995 = n34994 ^ n34474 ;
  assign n34996 = ~n34991 & n34995 ;
  assign n34997 = n34996 ^ n34990 ;
  assign n34988 = n34732 ^ n34731 ;
  assign n34989 = n34988 ^ n34560 ;
  assign n35147 = n34997 ^ n34989 ;
  assign n35148 = n33704 & n35147 ;
  assign n35149 = n35148 ^ n34560 ;
  assign n35200 = n35149 ^ n33397 ;
  assign n35029 = n35028 ^ n33399 ;
  assign n35144 = n35143 ^ n35028 ;
  assign n35145 = n35029 & ~n35144 ;
  assign n35146 = n35145 ^ n33399 ;
  assign n35201 = n35200 ^ n35146 ;
  assign n35202 = n35201 ^ x351 ;
  assign n35321 = n35296 ^ n35202 ;
  assign n35422 = n35358 ^ n35321 ;
  assign n35570 = n35422 ^ n35055 ;
  assign n35390 = n35389 ^ n34885 ;
  assign n35419 = n35418 ^ n35389 ;
  assign n35420 = n35390 & ~n35419 ;
  assign n35421 = n35420 ^ n34885 ;
  assign n35571 = n35570 ^ n35421 ;
  assign n35572 = ~n34222 & n35571 ;
  assign n35573 = n35572 ^ n35055 ;
  assign n35574 = n35573 ^ n33339 ;
  assign n35714 = n35621 ^ n35574 ;
  assign n35715 = n35714 ^ x32 ;
  assign n35865 = n35747 ^ n35715 ;
  assign n35866 = n35864 & ~n35865 ;
  assign n35748 = n35747 ^ n35714 ;
  assign n35749 = n35715 & ~n35748 ;
  assign n35750 = n35749 ^ x32 ;
  assign n35867 = n35750 ^ x47 ;
  assign n35622 = n35621 ^ n35573 ;
  assign n35623 = ~n35574 & n35622 ;
  assign n35624 = n35623 ^ n33339 ;
  assign n35712 = n35624 ^ n33336 ;
  assign n35423 = n35422 ^ n35421 ;
  assign n35359 = n35321 & n35358 ;
  assign n35150 = n35149 ^ n35146 ;
  assign n34987 = n34735 ^ n34733 ;
  assign n35021 = n34987 ^ n34470 ;
  assign n34998 = n34997 ^ n34988 ;
  assign n34999 = n34989 & ~n34998 ;
  assign n35000 = n34999 ^ n34560 ;
  assign n35022 = n35021 ^ n35000 ;
  assign n35023 = ~n33700 & ~n35022 ;
  assign n35024 = n35023 ^ n34470 ;
  assign n35151 = n35024 ^ n33397 ;
  assign n35152 = n35151 ^ n35146 ;
  assign n35153 = n35152 ^ n35024 ;
  assign n35154 = n35150 & ~n35153 ;
  assign n35155 = n35154 ^ n35151 ;
  assign n35199 = n35155 ^ n33393 ;
  assign n35319 = n35199 ^ x350 ;
  assign n35297 = n35296 ^ n35201 ;
  assign n35298 = ~n35202 & n35297 ;
  assign n35299 = n35298 ^ x351 ;
  assign n35320 = n35319 ^ n35299 ;
  assign n35424 = n35359 ^ n35320 ;
  assign n35425 = n35424 ^ n35055 ;
  assign n35426 = n35425 ^ n35421 ;
  assign n35427 = n35426 ^ n35424 ;
  assign n35428 = ~n35423 & n35427 ;
  assign n35429 = n35428 ^ n35425 ;
  assign n35566 = n35429 ^ n35065 ;
  assign n35567 = n34229 & n35566 ;
  assign n35568 = n35567 ^ n35065 ;
  assign n35713 = n35712 ^ n35568 ;
  assign n35868 = n35867 ^ n35713 ;
  assign n35869 = n35866 & ~n35868 ;
  assign n35751 = n35750 ^ n35713 ;
  assign n35754 = n35713 ^ x47 ;
  assign n35755 = ~n35751 & n35754 ;
  assign n35360 = n35320 & n35359 ;
  assign n35300 = n35299 ^ n35199 ;
  assign n35301 = n35299 ^ x350 ;
  assign n35302 = n35300 & n35301 ;
  assign n35303 = n35302 ^ x350 ;
  assign n35001 = n35000 ^ n34987 ;
  assign n35002 = n34737 ^ n34736 ;
  assign n35003 = n35002 ^ n34470 ;
  assign n35004 = n35003 ^ n34987 ;
  assign n35005 = n35004 ^ n35002 ;
  assign n35006 = n35001 & ~n35005 ;
  assign n35007 = n35006 ^ n35003 ;
  assign n35018 = n35007 ^ n34466 ;
  assign n35019 = ~n33696 & ~n35018 ;
  assign n35020 = n35019 ^ n34466 ;
  assign n35196 = n35020 ^ n33390 ;
  assign n35025 = n35024 ^ n33393 ;
  assign n35156 = ~n35025 & ~n35155 ;
  assign n35157 = n35156 ^ n33393 ;
  assign n35197 = n35196 ^ n35157 ;
  assign n35198 = n35197 ^ x349 ;
  assign n35318 = n35303 ^ n35198 ;
  assign n35430 = n35360 ^ n35318 ;
  assign n35432 = n35430 ^ n35065 ;
  assign n35431 = n35430 ^ n35424 ;
  assign n35433 = n35432 ^ n35431 ;
  assign n35434 = ~n35429 & n35433 ;
  assign n35435 = n35434 ^ n35432 ;
  assign n35629 = n35435 ^ n35051 ;
  assign n35630 = n34168 & ~n35629 ;
  assign n35631 = n35630 ^ n35051 ;
  assign n35569 = n35568 ^ n33336 ;
  assign n35625 = n35624 ^ n35568 ;
  assign n35626 = ~n35569 & n35625 ;
  assign n35627 = n35626 ^ n33336 ;
  assign n35628 = n35627 ^ n33760 ;
  assign n35710 = n35631 ^ n35628 ;
  assign n35752 = n35710 ^ x47 ;
  assign n35756 = n35755 ^ n35752 ;
  assign n35870 = n35756 ^ x46 ;
  assign n35871 = ~n35869 & ~n35870 ;
  assign n35361 = ~n35318 & n35360 ;
  assign n35158 = n35157 ^ n35020 ;
  assign n35008 = n34740 ^ n34738 ;
  assign n35010 = n35008 ^ n34466 ;
  assign n35009 = n35008 ^ n35002 ;
  assign n35011 = n35010 ^ n35009 ;
  assign n35012 = n35007 & ~n35011 ;
  assign n35013 = n35012 ^ n35010 ;
  assign n35014 = n35013 ^ n34575 ;
  assign n35015 = ~n33692 & n35014 ;
  assign n35016 = n35015 ^ n34575 ;
  assign n35159 = n35016 ^ n33390 ;
  assign n35160 = n35159 ^ n35020 ;
  assign n35161 = n35160 ^ n35016 ;
  assign n35162 = n35158 & ~n35161 ;
  assign n35163 = n35162 ^ n35159 ;
  assign n35195 = n35163 ^ n33387 ;
  assign n35316 = n35195 ^ x348 ;
  assign n35304 = n35303 ^ n35197 ;
  assign n35305 = n35198 & ~n35304 ;
  assign n35306 = n35305 ^ x349 ;
  assign n35317 = n35316 ^ n35306 ;
  assign n35436 = n35361 ^ n35317 ;
  assign n35438 = n35436 ^ n35051 ;
  assign n35437 = n35436 ^ n35430 ;
  assign n35439 = n35438 ^ n35437 ;
  assign n35440 = n35435 & ~n35439 ;
  assign n35441 = n35440 ^ n35438 ;
  assign n35636 = n35441 ^ n35047 ;
  assign n35637 = ~n34245 & ~n35636 ;
  assign n35638 = n35637 ^ n35047 ;
  assign n35632 = n35631 ^ n35627 ;
  assign n35633 = ~n35628 & n35632 ;
  assign n35634 = n35633 ^ n33760 ;
  assign n35635 = n35634 ^ n33805 ;
  assign n35760 = n35638 ^ n35635 ;
  assign n35711 = n35710 ^ x46 ;
  assign n35757 = ~n35711 & n35756 ;
  assign n35758 = n35757 ^ x46 ;
  assign n35759 = n35758 ^ x45 ;
  assign n35872 = n35760 ^ n35759 ;
  assign n35873 = ~n35871 & n35872 ;
  assign n35362 = n35317 & n35361 ;
  assign n35307 = n35306 ^ n35195 ;
  assign n35308 = n35306 ^ x348 ;
  assign n35309 = n35307 & n35308 ;
  assign n35310 = n35309 ^ x348 ;
  assign n35168 = n35008 ^ n34575 ;
  assign n35169 = ~n35013 & n35168 ;
  assign n35170 = n35169 ^ n34575 ;
  assign n35166 = n34742 ^ n34741 ;
  assign n35167 = n35166 ^ n34463 ;
  assign n35171 = n35170 ^ n35167 ;
  assign n35172 = n33871 & n35171 ;
  assign n35173 = n35172 ^ n34463 ;
  assign n35192 = n35173 ^ n33462 ;
  assign n35017 = n35016 ^ n33387 ;
  assign n35164 = n35017 & n35163 ;
  assign n35165 = n35164 ^ n33387 ;
  assign n35193 = n35192 ^ n35165 ;
  assign n35194 = n35193 ^ x347 ;
  assign n35315 = n35310 ^ n35194 ;
  assign n35387 = n35362 ^ n35315 ;
  assign n35443 = n35387 ^ n35047 ;
  assign n35442 = n35436 ^ n35387 ;
  assign n35444 = n35443 ^ n35442 ;
  assign n35445 = ~n35441 & ~n35444 ;
  assign n35446 = n35445 ^ n35443 ;
  assign n35563 = n35446 ^ n35080 ;
  assign n35564 = ~n34320 & n35563 ;
  assign n35565 = n35564 ^ n35080 ;
  assign n35708 = n35565 ^ n33756 ;
  assign n35639 = n35638 ^ n35634 ;
  assign n35640 = n35635 & n35639 ;
  assign n35641 = n35640 ^ n33805 ;
  assign n35709 = n35708 ^ n35641 ;
  assign n35850 = n35709 ^ x44 ;
  assign n35761 = n35760 ^ n35758 ;
  assign n35762 = n35759 & n35761 ;
  assign n35763 = n35762 ^ x45 ;
  assign n35851 = n35850 ^ n35763 ;
  assign n36015 = n35873 ^ n35851 ;
  assign n36209 = n36015 ^ n35509 ;
  assign n36016 = n35509 & ~n36015 ;
  assign n35874 = n35851 & n35873 ;
  assign n35764 = n35763 ^ n35709 ;
  assign n35765 = n35763 ^ x44 ;
  assign n35766 = n35764 & n35765 ;
  assign n35767 = n35766 ^ x44 ;
  assign n35642 = n35641 ^ n35565 ;
  assign n35643 = n35641 ^ n33756 ;
  assign n35644 = n35642 & n35643 ;
  assign n35645 = n35644 ^ n33756 ;
  assign n35705 = n35645 ^ n33752 ;
  assign n35363 = n35315 & n35362 ;
  assign n35311 = n35310 ^ n35193 ;
  assign n35312 = ~n35194 & n35311 ;
  assign n35313 = n35312 ^ x347 ;
  assign n35174 = n35173 ^ n35165 ;
  assign n35181 = n34745 ^ n34743 ;
  assign n35175 = n35170 ^ n35166 ;
  assign n35176 = n34592 ^ n34463 ;
  assign n35177 = n35176 ^ n34592 ;
  assign n35178 = n35177 ^ n35166 ;
  assign n35179 = ~n35175 & n35178 ;
  assign n35180 = n35179 ^ n35176 ;
  assign n35182 = n35181 ^ n35180 ;
  assign n35183 = n33688 & n35182 ;
  assign n35184 = n35183 ^ n34592 ;
  assign n35185 = n35184 ^ n33462 ;
  assign n35186 = n35185 ^ n35165 ;
  assign n35187 = n35186 ^ n35184 ;
  assign n35188 = ~n35174 & ~n35187 ;
  assign n35189 = n35188 ^ n35185 ;
  assign n35190 = n35189 ^ n33475 ;
  assign n35191 = n35190 ^ x346 ;
  assign n35314 = n35313 ^ n35191 ;
  assign n35449 = n35363 ^ n35314 ;
  assign n35558 = n35449 ^ n35043 ;
  assign n35388 = n35387 ^ n35080 ;
  assign n35447 = ~n35388 & n35446 ;
  assign n35448 = n35447 ^ n35080 ;
  assign n35559 = n35558 ^ n35448 ;
  assign n35560 = n34506 & n35559 ;
  assign n35561 = n35560 ^ n35043 ;
  assign n35706 = n35705 ^ n35561 ;
  assign n35707 = n35706 ^ x43 ;
  assign n35849 = n35767 ^ n35707 ;
  assign n36014 = n35874 ^ n35849 ;
  assign n36017 = n36016 ^ n36014 ;
  assign n35875 = ~n35849 & n35874 ;
  assign n35450 = n35449 ^ n35448 ;
  assign n35379 = n35184 ^ n33475 ;
  assign n35380 = n35189 & ~n35379 ;
  assign n35381 = n35380 ^ n33475 ;
  assign n35374 = n34747 ^ n34746 ;
  assign n35370 = n34712 ^ n34592 ;
  assign n35369 = n35181 ^ n34712 ;
  assign n35371 = n35370 ^ n35369 ;
  assign n35372 = n35180 & n35371 ;
  assign n35373 = n35372 ^ n35370 ;
  assign n35375 = n35374 ^ n35373 ;
  assign n35376 = ~n33887 & ~n35375 ;
  assign n35377 = n35376 ^ n34712 ;
  assign n35378 = n35377 ^ n33542 ;
  assign n35382 = n35381 ^ n35378 ;
  assign n35383 = n35382 ^ x345 ;
  assign n35365 = n35313 ^ n35190 ;
  assign n35366 = n35313 ^ x346 ;
  assign n35367 = ~n35365 & n35366 ;
  assign n35368 = n35367 ^ x346 ;
  assign n35384 = n35383 ^ n35368 ;
  assign n35364 = ~n35314 & n35363 ;
  assign n35385 = n35384 ^ n35364 ;
  assign n35451 = n35385 ^ n35043 ;
  assign n35452 = n35451 ^ n35448 ;
  assign n35453 = n35452 ^ n35385 ;
  assign n35454 = ~n35450 & ~n35453 ;
  assign n35455 = n35454 ^ n35451 ;
  assign n35555 = n35455 ^ n35091 ;
  assign n35556 = n34420 & n35555 ;
  assign n35557 = n35556 ^ n35091 ;
  assign n35771 = n35557 ^ n33749 ;
  assign n35562 = n35561 ^ n33752 ;
  assign n35646 = n35645 ^ n35561 ;
  assign n35647 = n35562 & ~n35646 ;
  assign n35648 = n35647 ^ n33752 ;
  assign n35772 = n35771 ^ n35648 ;
  assign n35847 = n35772 ^ x42 ;
  assign n35768 = n35767 ^ n35706 ;
  assign n35769 = n35707 & ~n35768 ;
  assign n35770 = n35769 ^ x43 ;
  assign n35848 = n35847 ^ n35770 ;
  assign n36012 = n35875 ^ n35848 ;
  assign n36018 = n36012 ^ n35591 ;
  assign n36019 = n36018 ^ n36014 ;
  assign n36020 = n36019 ^ n36012 ;
  assign n36021 = ~n36017 & ~n36020 ;
  assign n36022 = n36021 ^ n36018 ;
  assign n36205 = n36022 ^ n35600 ;
  assign n36206 = ~n34900 & ~n36205 ;
  assign n36207 = n36206 ^ n35600 ;
  assign n36208 = n36207 ^ n34185 ;
  assign n36213 = n36016 ^ n35591 ;
  assign n36214 = n36213 ^ n36014 ;
  assign n36215 = n34909 & n36214 ;
  assign n36216 = n36215 ^ n35591 ;
  assign n36210 = ~n34904 & n36209 ;
  assign n36211 = n36210 ^ n35509 ;
  assign n36212 = ~n34188 & ~n36211 ;
  assign n36217 = n36216 ^ n36212 ;
  assign n36218 = n36216 ^ n34193 ;
  assign n36219 = ~n36217 & n36218 ;
  assign n36220 = n36219 ^ n34193 ;
  assign n36221 = n36220 ^ n36207 ;
  assign n36222 = ~n36208 & n36221 ;
  assign n36223 = n36222 ^ n34185 ;
  assign n36224 = n36223 ^ n35408 ;
  assign n36013 = n36012 ^ n35600 ;
  assign n36023 = ~n36013 & ~n36022 ;
  assign n36024 = n36023 ^ n35600 ;
  assign n36202 = n36024 ^ n35585 ;
  assign n35876 = n35848 & ~n35875 ;
  assign n35773 = n35772 ^ n35770 ;
  assign n35649 = n35648 ^ n35557 ;
  assign n35650 = n35648 ^ n33749 ;
  assign n35651 = ~n35649 & n35650 ;
  assign n35652 = n35651 ^ n33749 ;
  assign n35702 = n35652 ^ n33823 ;
  assign n35474 = n35382 ^ n35364 ;
  assign n35477 = n35474 ^ n35368 ;
  assign n35478 = x345 & ~n35477 ;
  assign n35475 = n35368 ^ n35364 ;
  assign n35476 = ~n35474 & n35475 ;
  assign n35479 = n35478 ^ n35476 ;
  assign n35470 = n34778 ^ n33581 ;
  assign n35469 = n33542 ^ x344 ;
  assign n35471 = n35470 ^ n35469 ;
  assign n35464 = n34778 ^ n34748 ;
  assign n35465 = n35464 ^ n34749 ;
  assign n35466 = n35465 ^ n35374 ;
  assign n35462 = n35374 ^ n34712 ;
  assign n35463 = n35373 & ~n35462 ;
  assign n35467 = n35466 ^ n35463 ;
  assign n35468 = ~n33903 & ~n35467 ;
  assign n35472 = n35471 ^ n35468 ;
  assign n35459 = n35381 ^ n35377 ;
  assign n35460 = n35381 ^ n33542 ;
  assign n35461 = ~n35459 & n35460 ;
  assign n35473 = n35472 ^ n35461 ;
  assign n35480 = n35479 ^ n35473 ;
  assign n35386 = n35385 ^ n35091 ;
  assign n35456 = n35386 & ~n35455 ;
  assign n35457 = n35456 ^ n35091 ;
  assign n35458 = n35457 ^ n35097 ;
  assign n35653 = n35480 ^ n35458 ;
  assign n35654 = ~n34416 & ~n35653 ;
  assign n35655 = n35654 ^ n35097 ;
  assign n35703 = n35702 ^ n35655 ;
  assign n35774 = n35703 ^ x42 ;
  assign n35775 = n35774 ^ n35770 ;
  assign n35776 = n35775 ^ n35703 ;
  assign n35777 = ~n35773 & n35776 ;
  assign n35778 = n35777 ^ n35774 ;
  assign n35846 = n35778 ^ x41 ;
  assign n36025 = n35876 ^ n35846 ;
  assign n36203 = n36202 ^ n36025 ;
  assign n36204 = ~n34896 & n36203 ;
  assign n36225 = n36224 ^ n36204 ;
  assign n36226 = n36223 ^ n34204 ;
  assign n36227 = ~n36225 & ~n36226 ;
  assign n36228 = n36227 ^ n34204 ;
  assign n36395 = n36228 ^ n34180 ;
  assign n35877 = n35846 & ~n35876 ;
  assign n35656 = n35655 ^ n35652 ;
  assign n35481 = n35480 ^ n35457 ;
  assign n35482 = n35458 & n35481 ;
  assign n35483 = n35482 ^ n35097 ;
  assign n35484 = n35483 ^ n34963 ;
  assign n35551 = n35484 ^ n35038 ;
  assign n35552 = n34413 & ~n35551 ;
  assign n35553 = n35552 ^ n35038 ;
  assign n35657 = n35553 ^ n33823 ;
  assign n35658 = n35657 ^ n35553 ;
  assign n35659 = n35658 ^ n35652 ;
  assign n35660 = ~n35656 & ~n35659 ;
  assign n35661 = n35660 ^ n35657 ;
  assign n35781 = n35661 ^ n33744 ;
  assign n35844 = n35781 ^ x40 ;
  assign n35704 = n35703 ^ x41 ;
  assign n35779 = ~n35704 & n35778 ;
  assign n35780 = n35779 ^ x41 ;
  assign n35845 = n35844 ^ n35780 ;
  assign n36030 = n35877 ^ n35845 ;
  assign n36229 = n36030 ^ n35609 ;
  assign n36026 = n36025 ^ n36024 ;
  assign n36027 = n36025 ^ n35585 ;
  assign n36028 = ~n36026 & n36027 ;
  assign n36029 = n36028 ^ n35585 ;
  assign n36230 = n36229 ^ n36029 ;
  assign n36231 = ~n34892 & n36230 ;
  assign n36232 = n36231 ^ n35609 ;
  assign n36396 = n36395 ^ n36232 ;
  assign n36397 = n36396 ^ x259 ;
  assign n36399 = n35395 ^ n34797 ;
  assign n36400 = n36399 ^ n36210 ;
  assign n36401 = x263 & n36400 ;
  assign n36402 = n36401 ^ x262 ;
  assign n36403 = n36212 ^ n34193 ;
  assign n36404 = n36403 ^ n36216 ;
  assign n36405 = n36404 ^ n36401 ;
  assign n36406 = n36402 & ~n36405 ;
  assign n36407 = n36406 ^ x262 ;
  assign n36398 = n36220 ^ n36208 ;
  assign n36408 = n36407 ^ n36398 ;
  assign n36409 = n36225 ^ n34204 ;
  assign n36410 = n36409 ^ x261 ;
  assign n36411 = n36410 ^ n36398 ;
  assign n36412 = n36411 ^ n36409 ;
  assign n36413 = n36408 & ~n36412 ;
  assign n36414 = n36413 ^ n36410 ;
  assign n36416 = n36396 ^ x260 ;
  assign n36415 = n36409 ^ n36396 ;
  assign n36417 = n36416 ^ n36415 ;
  assign n36418 = n36414 & ~n36417 ;
  assign n36419 = n36418 ^ n36416 ;
  assign n36420 = n36397 & ~n36419 ;
  assign n36421 = n36420 ^ x259 ;
  assign n36422 = n36421 ^ x258 ;
  assign n36031 = n36030 ^ n36029 ;
  assign n35782 = n35781 ^ n35780 ;
  assign n35554 = n35553 ^ n33744 ;
  assign n35662 = ~n35554 & ~n35661 ;
  assign n35663 = n35662 ^ n33744 ;
  assign n35488 = n34964 ^ n34963 ;
  assign n35546 = n35488 ^ n35107 ;
  assign n35485 = n35038 ^ n34963 ;
  assign n35486 = ~n35484 & ~n35485 ;
  assign n35487 = n35486 ^ n35038 ;
  assign n35547 = n35546 ^ n35487 ;
  assign n35548 = ~n34409 & n35547 ;
  assign n35549 = n35548 ^ n35107 ;
  assign n35550 = n35549 ^ n33740 ;
  assign n35783 = n35663 ^ n35550 ;
  assign n35784 = n35783 ^ x40 ;
  assign n35785 = n35784 ^ n35780 ;
  assign n35786 = n35785 ^ n35783 ;
  assign n35787 = ~n35782 & n35786 ;
  assign n35788 = n35787 ^ n35784 ;
  assign n35879 = n35788 ^ x55 ;
  assign n35878 = n35845 & ~n35877 ;
  assign n36010 = n35879 ^ n35878 ;
  assign n36032 = n36010 ^ n35609 ;
  assign n36033 = n36032 ^ n36010 ;
  assign n36034 = n36033 ^ n36029 ;
  assign n36035 = n36031 & n36034 ;
  assign n36036 = n36035 ^ n36032 ;
  assign n36237 = n36036 ^ n35581 ;
  assign n36238 = ~n34888 & ~n36237 ;
  assign n36239 = n36238 ^ n35581 ;
  assign n36241 = n36239 ^ n34176 ;
  assign n36233 = n36232 ^ n36228 ;
  assign n36234 = n36232 ^ n34180 ;
  assign n36235 = ~n36233 & ~n36234 ;
  assign n36236 = n36235 ^ n34180 ;
  assign n36423 = n36241 ^ n36236 ;
  assign n36424 = n36423 ^ n36421 ;
  assign n36425 = n36422 & ~n36424 ;
  assign n36426 = n36425 ^ x258 ;
  assign n35664 = n35663 ^ n35549 ;
  assign n35665 = n35550 & ~n35664 ;
  assign n35666 = n35665 ^ n33740 ;
  assign n35489 = n35488 ^ n35487 ;
  assign n35492 = n35487 ^ n35107 ;
  assign n35493 = ~n35489 & ~n35492 ;
  assign n34984 = n34966 ^ n34965 ;
  assign n35490 = n35107 ^ n34984 ;
  assign n35494 = n35493 ^ n35490 ;
  assign n35542 = n35494 ^ n34985 ;
  assign n35543 = n34406 & ~n35542 ;
  assign n35544 = n35543 ^ n34985 ;
  assign n35545 = n35544 ^ n33735 ;
  assign n35789 = n35666 ^ n35545 ;
  assign n35791 = n35789 ^ x55 ;
  assign n35790 = n35789 ^ n35783 ;
  assign n35792 = n35791 ^ n35790 ;
  assign n35793 = ~n35788 & n35792 ;
  assign n35794 = n35793 ^ n35791 ;
  assign n35881 = n35794 ^ x54 ;
  assign n35880 = n35878 & n35879 ;
  assign n36009 = n35881 ^ n35880 ;
  assign n36244 = n36009 ^ n35576 ;
  assign n36011 = n36010 ^ n35581 ;
  assign n36037 = n36011 & ~n36036 ;
  assign n36038 = n36037 ^ n35581 ;
  assign n36245 = n36244 ^ n36038 ;
  assign n36246 = ~n34885 & ~n36245 ;
  assign n36247 = n36246 ^ n35576 ;
  assign n36393 = n36247 ^ n34172 ;
  assign n36240 = n36239 ^ n36236 ;
  assign n36242 = n36240 & n36241 ;
  assign n36243 = n36242 ^ n34176 ;
  assign n36394 = n36393 ^ n36243 ;
  assign n36427 = n36426 ^ n36394 ;
  assign n36248 = n36247 ^ n36243 ;
  assign n36039 = n36038 ^ n36009 ;
  assign n36040 = n36038 ^ n35576 ;
  assign n36041 = n36039 & ~n36040 ;
  assign n36042 = n36041 ^ n35576 ;
  assign n35667 = n35666 ^ n35544 ;
  assign n35668 = ~n35545 & n35667 ;
  assign n35669 = n35668 ^ n33735 ;
  assign n35699 = n35669 ^ n33731 ;
  assign n34986 = n34985 ^ n34984 ;
  assign n35495 = ~n34986 & ~n35494 ;
  assign n35496 = n35495 ^ n34985 ;
  assign n34981 = n34969 ^ n34967 ;
  assign n34983 = n34982 ^ n34981 ;
  assign n35538 = n35496 ^ n34983 ;
  assign n35539 = n34403 & ~n35538 ;
  assign n35540 = n35539 ^ n34982 ;
  assign n35700 = n35699 ^ n35540 ;
  assign n35796 = n35700 ^ x54 ;
  assign n35795 = n35789 ^ n35700 ;
  assign n35797 = n35796 ^ n35795 ;
  assign n35798 = n35794 & ~n35797 ;
  assign n35799 = n35798 ^ n35796 ;
  assign n35883 = n35799 ^ x53 ;
  assign n35882 = n35880 & ~n35881 ;
  assign n36007 = n35883 ^ n35882 ;
  assign n36008 = n36007 ^ n35571 ;
  assign n36198 = n36042 ^ n36008 ;
  assign n36199 = ~n35055 & n36198 ;
  assign n36200 = n36199 ^ n35571 ;
  assign n36249 = n36200 ^ n34172 ;
  assign n36250 = n36249 ^ n36200 ;
  assign n36251 = n36250 ^ n36243 ;
  assign n36252 = n36248 & n36251 ;
  assign n36253 = n36252 ^ n36249 ;
  assign n36391 = n36253 ^ n34222 ;
  assign n36428 = n36391 ^ x257 ;
  assign n36429 = n36428 ^ n36391 ;
  assign n36430 = n36429 ^ n36394 ;
  assign n36431 = ~n36427 & n36430 ;
  assign n36432 = n36431 ^ n36428 ;
  assign n36515 = n36432 ^ x256 ;
  assign n36516 = n36419 ^ x259 ;
  assign n36517 = n36400 ^ x263 ;
  assign n36518 = n36404 ^ x262 ;
  assign n36519 = n36518 ^ n36401 ;
  assign n36520 = ~n36517 & ~n36519 ;
  assign n36521 = n36407 ^ x261 ;
  assign n36522 = n36521 ^ n36398 ;
  assign n36523 = n36520 & n36522 ;
  assign n36524 = n36414 ^ x260 ;
  assign n36525 = n36523 & n36524 ;
  assign n36526 = n36516 & ~n36525 ;
  assign n36527 = n36423 ^ n36422 ;
  assign n36528 = n36526 & n36527 ;
  assign n36529 = n36394 ^ x257 ;
  assign n36530 = n36529 ^ n36426 ;
  assign n36531 = ~n36528 & ~n36530 ;
  assign n36532 = n36515 & ~n36531 ;
  assign n35541 = n35540 ^ n33731 ;
  assign n35670 = n35669 ^ n35540 ;
  assign n35671 = n35541 & ~n35670 ;
  assign n35672 = n35671 ^ n33731 ;
  assign n35697 = n35672 ^ n33727 ;
  assign n34980 = n34971 ^ n34970 ;
  assign n35533 = n35124 ^ n34980 ;
  assign n35497 = n35496 ^ n34981 ;
  assign n35498 = n34983 & n35497 ;
  assign n35499 = n35498 ^ n34982 ;
  assign n35534 = n35533 ^ n35499 ;
  assign n35535 = ~n34485 & n35534 ;
  assign n35536 = n35535 ^ n35124 ;
  assign n35698 = n35697 ^ n35536 ;
  assign n35885 = n35698 ^ x52 ;
  assign n35701 = n35700 ^ x53 ;
  assign n35800 = n35701 & ~n35799 ;
  assign n35801 = n35800 ^ x53 ;
  assign n35886 = n35885 ^ n35801 ;
  assign n35884 = ~n35882 & ~n35883 ;
  assign n36006 = n35886 ^ n35884 ;
  assign n36194 = n36006 ^ n35566 ;
  assign n36043 = n36042 ^ n36007 ;
  assign n36044 = n36008 & ~n36043 ;
  assign n36045 = n36044 ^ n35571 ;
  assign n36195 = n36194 ^ n36045 ;
  assign n36196 = ~n35065 & ~n36195 ;
  assign n36197 = n36196 ^ n35566 ;
  assign n36389 = n36197 ^ n34229 ;
  assign n36201 = n36200 ^ n34222 ;
  assign n36254 = ~n36201 & n36253 ;
  assign n36255 = n36254 ^ n34222 ;
  assign n36390 = n36389 ^ n36255 ;
  assign n36533 = n36390 ^ x271 ;
  assign n36392 = n36391 ^ x256 ;
  assign n36433 = n36392 & ~n36432 ;
  assign n36434 = n36433 ^ x256 ;
  assign n36534 = n36533 ^ n36434 ;
  assign n36535 = n36532 & ~n36534 ;
  assign n36435 = n36434 ^ n36390 ;
  assign n36436 = n36434 ^ x271 ;
  assign n36437 = n36435 & n36436 ;
  assign n36438 = n36437 ^ x271 ;
  assign n36256 = n36255 ^ n36197 ;
  assign n36257 = n36255 ^ n34229 ;
  assign n36258 = n36256 & ~n36257 ;
  assign n36259 = n36258 ^ n34229 ;
  assign n35887 = ~n35884 & ~n35886 ;
  assign n35500 = n35499 ^ n34980 ;
  assign n34977 = n34972 ^ n34962 ;
  assign n35501 = n35124 ^ n34977 ;
  assign n35502 = n35501 ^ n34980 ;
  assign n35503 = n35502 ^ n34977 ;
  assign n35504 = ~n35500 & n35503 ;
  assign n35505 = n35504 ^ n35501 ;
  assign n35677 = n35505 ^ n34978 ;
  assign n35678 = ~n34543 & ~n35677 ;
  assign n35679 = n35678 ^ n34978 ;
  assign n35537 = n35536 ^ n33727 ;
  assign n35673 = n35672 ^ n35536 ;
  assign n35674 = ~n35537 & ~n35673 ;
  assign n35675 = n35674 ^ n33727 ;
  assign n35676 = n35675 ^ n33722 ;
  assign n35806 = n35679 ^ n35676 ;
  assign n35842 = n35806 ^ x51 ;
  assign n35802 = n35801 ^ n35698 ;
  assign n35803 = n35801 ^ x52 ;
  assign n35804 = n35802 & n35803 ;
  assign n35805 = n35804 ^ x52 ;
  assign n35843 = n35842 ^ n35805 ;
  assign n36050 = n35887 ^ n35843 ;
  assign n36189 = n36050 ^ n35629 ;
  assign n36046 = n36045 ^ n36006 ;
  assign n36047 = n36045 ^ n35566 ;
  assign n36048 = n36046 & n36047 ;
  assign n36049 = n36048 ^ n35566 ;
  assign n36190 = n36189 ^ n36049 ;
  assign n36191 = ~n35051 & n36190 ;
  assign n36192 = n36191 ^ n35629 ;
  assign n36193 = n36192 ^ n34168 ;
  assign n36387 = n36259 ^ n36193 ;
  assign n36388 = n36387 ^ x270 ;
  assign n36536 = n36438 ^ n36388 ;
  assign n36537 = ~n36535 & n36536 ;
  assign n36051 = n36050 ^ n36049 ;
  assign n35888 = n35843 & n35887 ;
  assign n35807 = n35806 ^ n35805 ;
  assign n35811 = n35805 ^ x51 ;
  assign n35812 = ~n35807 & n35811 ;
  assign n34979 = n34978 ^ n34977 ;
  assign n35506 = ~n34979 & ~n35505 ;
  assign n35507 = n35506 ^ n34978 ;
  assign n34974 = n34973 ^ n34961 ;
  assign n34976 = n34975 ^ n34974 ;
  assign n35508 = n35507 ^ n34976 ;
  assign n35684 = n34401 & n35508 ;
  assign n35685 = n35684 ^ n34975 ;
  assign n35680 = n35679 ^ n35675 ;
  assign n35681 = ~n35676 & ~n35680 ;
  assign n35682 = n35681 ^ n33722 ;
  assign n35683 = n35682 ^ n33717 ;
  assign n35808 = n35685 ^ n35683 ;
  assign n35809 = n35808 ^ x51 ;
  assign n35813 = n35812 ^ n35809 ;
  assign n35841 = n35813 ^ x50 ;
  assign n36052 = n35888 ^ n35841 ;
  assign n36053 = n36052 ^ n35629 ;
  assign n36054 = n36053 ^ n36052 ;
  assign n36055 = n36054 ^ n36049 ;
  assign n36056 = n36051 & ~n36055 ;
  assign n36057 = n36056 ^ n36053 ;
  assign n36186 = n36057 ^ n35636 ;
  assign n36187 = n35047 & ~n36186 ;
  assign n36188 = n36187 ^ n35636 ;
  assign n36385 = n36188 ^ n34245 ;
  assign n36260 = n36259 ^ n36192 ;
  assign n36261 = ~n36193 & n36260 ;
  assign n36262 = n36261 ^ n34168 ;
  assign n36386 = n36385 ^ n36262 ;
  assign n36538 = n36386 ^ x269 ;
  assign n36439 = n36438 ^ n36387 ;
  assign n36440 = ~n36388 & n36439 ;
  assign n36441 = n36440 ^ x270 ;
  assign n36539 = n36538 ^ n36441 ;
  assign n36540 = n36537 & ~n36539 ;
  assign n36442 = n36441 ^ n36386 ;
  assign n36443 = n36441 ^ x269 ;
  assign n36444 = ~n36442 & n36443 ;
  assign n36445 = n36444 ^ x269 ;
  assign n36541 = n36445 ^ x268 ;
  assign n36263 = n36262 ^ n36188 ;
  assign n36264 = n36262 ^ n34245 ;
  assign n36265 = n36263 & ~n36264 ;
  assign n36266 = n36265 ^ n34245 ;
  assign n35686 = n35685 ^ n35682 ;
  assign n35687 = ~n35683 & n35686 ;
  assign n35688 = n35687 ^ n33717 ;
  assign n35694 = n35688 ^ n33712 ;
  assign n35521 = n35323 ^ n35322 ;
  assign n35517 = n34975 ^ n34884 ;
  assign n35514 = n35507 ^ n34974 ;
  assign n35515 = n35507 ^ n34975 ;
  assign n35516 = n35514 & n35515 ;
  assign n35518 = n35517 ^ n35516 ;
  assign n35529 = n35521 ^ n35518 ;
  assign n35530 = ~n34478 & n35529 ;
  assign n35531 = n35530 ^ n34884 ;
  assign n35695 = n35694 ^ n35531 ;
  assign n35815 = n35695 ^ x50 ;
  assign n35814 = n35808 ^ n35695 ;
  assign n35816 = n35815 ^ n35814 ;
  assign n35817 = ~n35813 & n35816 ;
  assign n35818 = n35817 ^ n35815 ;
  assign n35890 = n35818 ^ x49 ;
  assign n35889 = n35841 & n35888 ;
  assign n36004 = n35890 ^ n35889 ;
  assign n36059 = n36004 ^ n35636 ;
  assign n36058 = n36052 ^ n36004 ;
  assign n36060 = n36059 ^ n36058 ;
  assign n36061 = ~n36057 & n36060 ;
  assign n36062 = n36061 ^ n36059 ;
  assign n36182 = n36062 ^ n35563 ;
  assign n36183 = n35080 & n36182 ;
  assign n36184 = n36183 ^ n35563 ;
  assign n36185 = n36184 ^ n34320 ;
  assign n36383 = n36266 ^ n36185 ;
  assign n36542 = n36541 ^ n36383 ;
  assign n36543 = n36540 & ~n36542 ;
  assign n35532 = n35531 ^ n33712 ;
  assign n35689 = n35688 ^ n35531 ;
  assign n35690 = ~n35532 & ~n35689 ;
  assign n35691 = n35690 ^ n33712 ;
  assign n35692 = n35691 ^ n33708 ;
  assign n35519 = n35325 ^ n35324 ;
  assign n35520 = n35519 ^ n34884 ;
  assign n35522 = n35521 ^ n35520 ;
  assign n35523 = n35522 ^ n35519 ;
  assign n35524 = n35518 & ~n35523 ;
  assign n35525 = n35524 ^ n35520 ;
  assign n35526 = n35525 ^ n35026 ;
  assign n35527 = n34474 & n35526 ;
  assign n35528 = n35527 ^ n35026 ;
  assign n35693 = n35692 ^ n35528 ;
  assign n35892 = n35693 ^ x48 ;
  assign n35696 = n35695 ^ x49 ;
  assign n35819 = n35696 & ~n35818 ;
  assign n35820 = n35819 ^ x49 ;
  assign n35893 = n35892 ^ n35820 ;
  assign n35891 = n35889 & n35890 ;
  assign n36066 = n35893 ^ n35891 ;
  assign n36005 = n36004 ^ n35563 ;
  assign n36063 = ~n36005 & ~n36062 ;
  assign n36064 = n36063 ^ n35563 ;
  assign n36065 = n36064 ^ n35559 ;
  assign n36271 = n36066 ^ n36065 ;
  assign n36272 = ~n35043 & n36271 ;
  assign n36273 = n36272 ^ n35559 ;
  assign n36267 = n36266 ^ n36184 ;
  assign n36268 = ~n36185 & n36267 ;
  assign n36269 = n36268 ^ n34320 ;
  assign n36270 = n36269 ^ n34506 ;
  assign n36450 = n36273 ^ n36270 ;
  assign n36384 = n36383 ^ x268 ;
  assign n36446 = n36445 ^ n36383 ;
  assign n36447 = n36384 & ~n36446 ;
  assign n36448 = n36447 ^ x268 ;
  assign n36449 = n36448 ^ x267 ;
  assign n36544 = n36450 ^ n36449 ;
  assign n36545 = n36543 & n36544 ;
  assign n36067 = n36066 ^ n36064 ;
  assign n36068 = n36065 & ~n36067 ;
  assign n36069 = n36068 ^ n35559 ;
  assign n35894 = ~n35891 & ~n35893 ;
  assign n35821 = n35820 ^ n35693 ;
  assign n35831 = n35691 ^ n35528 ;
  assign n35832 = ~n35692 & n35831 ;
  assign n35833 = n35832 ^ n33708 ;
  assign n35825 = n35327 ^ n35326 ;
  assign n35826 = n35825 ^ n35147 ;
  assign n35822 = n35519 ^ n35026 ;
  assign n35823 = n35525 & ~n35822 ;
  assign n35824 = n35823 ^ n35026 ;
  assign n35827 = n35826 ^ n35824 ;
  assign n35828 = ~n34560 & n35827 ;
  assign n35829 = n35828 ^ n35147 ;
  assign n35830 = n35829 ^ n33704 ;
  assign n35834 = n35833 ^ n35830 ;
  assign n35835 = n35834 ^ x48 ;
  assign n35836 = n35835 ^ n35693 ;
  assign n35837 = n35836 ^ n35834 ;
  assign n35838 = ~n35821 & n35837 ;
  assign n35839 = n35838 ^ n35835 ;
  assign n35840 = n35839 ^ x63 ;
  assign n36002 = n35894 ^ n35840 ;
  assign n36003 = n36002 ^ n35555 ;
  assign n36179 = n36069 ^ n36003 ;
  assign n36180 = ~n35091 & n36179 ;
  assign n36181 = n36180 ^ n35555 ;
  assign n36381 = n36181 ^ n34420 ;
  assign n36274 = n36273 ^ n36269 ;
  assign n36275 = ~n36270 & n36274 ;
  assign n36276 = n36275 ^ n34506 ;
  assign n36382 = n36381 ^ n36276 ;
  assign n36546 = n36382 ^ x266 ;
  assign n36451 = n36450 ^ n36448 ;
  assign n36452 = n36449 & n36451 ;
  assign n36453 = n36452 ^ x267 ;
  assign n36547 = n36546 ^ n36453 ;
  assign n36548 = n36545 & ~n36547 ;
  assign n36454 = n36453 ^ n36382 ;
  assign n36455 = n36453 ^ x266 ;
  assign n36456 = ~n36454 & n36455 ;
  assign n36457 = n36456 ^ x266 ;
  assign n36549 = n36457 ^ x265 ;
  assign n36277 = n36276 ^ n36181 ;
  assign n36278 = n36276 ^ n34420 ;
  assign n36279 = ~n36277 & n36278 ;
  assign n36280 = n36279 ^ n34420 ;
  assign n35903 = n35329 ^ n35328 ;
  assign n35904 = n35903 ^ n35022 ;
  assign n35900 = n35825 ^ n35824 ;
  assign n35901 = ~n35826 & ~n35900 ;
  assign n35902 = n35901 ^ n35147 ;
  assign n35905 = n35904 ^ n35902 ;
  assign n35906 = ~n34470 & ~n35905 ;
  assign n35907 = n35906 ^ n35022 ;
  assign n35896 = n35833 ^ n35829 ;
  assign n35897 = n35830 & n35896 ;
  assign n35898 = n35897 ^ n33704 ;
  assign n35899 = n35898 ^ n33700 ;
  assign n35908 = n35907 ^ n35899 ;
  assign n35910 = n35908 ^ x63 ;
  assign n35909 = n35908 ^ n35834 ;
  assign n35911 = n35910 ^ n35909 ;
  assign n35912 = n35839 & ~n35911 ;
  assign n35913 = n35912 ^ n35910 ;
  assign n35914 = n35913 ^ x62 ;
  assign n35895 = n35840 & n35894 ;
  assign n36073 = n35914 ^ n35895 ;
  assign n36174 = n36073 ^ n35653 ;
  assign n36070 = n36069 ^ n36002 ;
  assign n36071 = n36003 & ~n36070 ;
  assign n36072 = n36071 ^ n35555 ;
  assign n36175 = n36174 ^ n36072 ;
  assign n36176 = ~n35097 & ~n36175 ;
  assign n36177 = n36176 ^ n35653 ;
  assign n36178 = n36177 ^ n34416 ;
  assign n36379 = n36280 ^ n36178 ;
  assign n36550 = n36549 ^ n36379 ;
  assign n36551 = n36548 & ~n36550 ;
  assign n36074 = n36073 ^ n36072 ;
  assign n35927 = n35332 ^ n35330 ;
  assign n35928 = n35927 ^ n35018 ;
  assign n35924 = n35903 ^ n35902 ;
  assign n35925 = ~n35904 & ~n35924 ;
  assign n35926 = n35925 ^ n35022 ;
  assign n35929 = n35928 ^ n35926 ;
  assign n35930 = ~n34466 & ~n35929 ;
  assign n35931 = n35930 ^ n35018 ;
  assign n35919 = n35907 ^ n33700 ;
  assign n35920 = n35907 ^ n35898 ;
  assign n35921 = n35919 & n35920 ;
  assign n35922 = n35921 ^ n33700 ;
  assign n35923 = n35922 ^ n33696 ;
  assign n35932 = n35931 ^ n35923 ;
  assign n35933 = n35932 ^ x61 ;
  assign n35916 = n35908 ^ x62 ;
  assign n35917 = ~n35913 & n35916 ;
  assign n35918 = n35917 ^ x62 ;
  assign n35934 = n35933 ^ n35918 ;
  assign n35915 = ~n35895 & n35914 ;
  assign n36000 = n35934 ^ n35915 ;
  assign n36075 = n36000 ^ n35653 ;
  assign n36076 = n36075 ^ n36000 ;
  assign n36077 = n36076 ^ n36072 ;
  assign n36078 = ~n36074 & ~n36077 ;
  assign n36079 = n36078 ^ n36075 ;
  assign n36171 = n36079 ^ n35551 ;
  assign n36172 = n35038 & ~n36171 ;
  assign n36173 = n36172 ^ n35551 ;
  assign n36377 = n36173 ^ n34413 ;
  assign n36281 = n36280 ^ n36177 ;
  assign n36282 = n36178 & n36281 ;
  assign n36283 = n36282 ^ n34416 ;
  assign n36378 = n36377 ^ n36283 ;
  assign n36552 = n36378 ^ x264 ;
  assign n36380 = n36379 ^ x265 ;
  assign n36458 = n36457 ^ n36379 ;
  assign n36459 = n36380 & ~n36458 ;
  assign n36460 = n36459 ^ x265 ;
  assign n36553 = n36552 ^ n36460 ;
  assign n36554 = ~n36551 & n36553 ;
  assign n36461 = n36460 ^ n36378 ;
  assign n36462 = n36460 ^ x264 ;
  assign n36463 = ~n36461 & n36462 ;
  assign n36464 = n36463 ^ x264 ;
  assign n36555 = n36464 ^ x279 ;
  assign n36001 = n36000 ^ n35551 ;
  assign n36080 = n36001 & ~n36079 ;
  assign n36081 = n36080 ^ n35551 ;
  assign n35945 = n35927 ^ n35926 ;
  assign n35946 = n35928 & ~n35945 ;
  assign n35947 = n35946 ^ n35018 ;
  assign n35943 = n35334 ^ n35333 ;
  assign n35944 = n35943 ^ n35014 ;
  assign n35948 = n35947 ^ n35944 ;
  assign n35949 = ~n34575 & n35948 ;
  assign n35950 = n35949 ^ n35014 ;
  assign n35951 = n35950 ^ n33692 ;
  assign n35939 = n35931 ^ n33696 ;
  assign n35940 = n35931 ^ n35922 ;
  assign n35941 = n35939 & ~n35940 ;
  assign n35942 = n35941 ^ n33696 ;
  assign n35952 = n35951 ^ n35942 ;
  assign n35953 = n35952 ^ x60 ;
  assign n35936 = n35932 ^ n35918 ;
  assign n35937 = ~n35933 & n35936 ;
  assign n35938 = n35937 ^ x61 ;
  assign n35954 = n35953 ^ n35938 ;
  assign n35935 = ~n35915 & n35934 ;
  assign n35998 = n35954 ^ n35935 ;
  assign n35999 = n35998 ^ n35547 ;
  assign n36288 = n36081 ^ n35999 ;
  assign n36289 = ~n35107 & ~n36288 ;
  assign n36290 = n36289 ^ n35547 ;
  assign n36374 = n36290 ^ n34409 ;
  assign n36284 = n36283 ^ n36173 ;
  assign n36285 = n36283 ^ n34413 ;
  assign n36286 = ~n36284 & ~n36285 ;
  assign n36287 = n36286 ^ n34413 ;
  assign n36375 = n36374 ^ n36287 ;
  assign n36556 = n36555 ^ n36375 ;
  assign n36557 = n36554 & ~n36556 ;
  assign n36291 = n36290 ^ n36287 ;
  assign n36082 = n36081 ^ n35998 ;
  assign n36083 = n35999 & n36082 ;
  assign n36084 = n36083 ^ n35547 ;
  assign n36166 = n36084 ^ n35542 ;
  assign n35969 = n35950 ^ n35942 ;
  assign n35970 = ~n35951 & n35969 ;
  assign n35971 = n35970 ^ n33692 ;
  assign n35963 = n35336 ^ n35335 ;
  assign n35964 = n35963 ^ n35171 ;
  assign n35959 = n35947 ^ n35943 ;
  assign n35960 = n35947 ^ n35014 ;
  assign n35961 = ~n35959 & ~n35960 ;
  assign n35962 = n35961 ^ n35014 ;
  assign n35965 = n35964 ^ n35962 ;
  assign n35966 = ~n34463 & ~n35965 ;
  assign n35967 = n35966 ^ n35171 ;
  assign n35968 = n35967 ^ n33871 ;
  assign n35972 = n35971 ^ n35968 ;
  assign n35973 = n35972 ^ x59 ;
  assign n35956 = n35952 ^ n35938 ;
  assign n35957 = n35953 & ~n35956 ;
  assign n35958 = n35957 ^ x60 ;
  assign n35974 = n35973 ^ n35958 ;
  assign n35955 = ~n35935 & n35954 ;
  assign n35996 = n35974 ^ n35955 ;
  assign n36167 = n36166 ^ n35996 ;
  assign n36168 = n34985 & ~n36167 ;
  assign n36169 = n36168 ^ n35542 ;
  assign n36292 = n36169 ^ n34409 ;
  assign n36293 = n36292 ^ n36169 ;
  assign n36294 = n36293 ^ n36287 ;
  assign n36295 = ~n36291 & ~n36294 ;
  assign n36296 = n36295 ^ n36292 ;
  assign n36373 = n36296 ^ n34406 ;
  assign n36558 = n36373 ^ x278 ;
  assign n36376 = n36375 ^ x279 ;
  assign n36465 = n36464 ^ n36375 ;
  assign n36466 = ~n36376 & n36465 ;
  assign n36467 = n36466 ^ x279 ;
  assign n36559 = n36558 ^ n36467 ;
  assign n36560 = n36557 & n36559 ;
  assign n36468 = n36467 ^ n36373 ;
  assign n36170 = n36169 ^ n34406 ;
  assign n36297 = ~n36170 & ~n36296 ;
  assign n36298 = n36297 ^ n34406 ;
  assign n36370 = n36298 ^ n34403 ;
  assign n35997 = n35996 ^ n35542 ;
  assign n36085 = n36084 ^ n35996 ;
  assign n36086 = ~n35997 & ~n36085 ;
  assign n36087 = n36086 ^ n35542 ;
  assign n35988 = n35971 ^ n35967 ;
  assign n35989 = n35968 & n35988 ;
  assign n35990 = n35989 ^ n33871 ;
  assign n35981 = n35963 ^ n35962 ;
  assign n35982 = ~n35964 & n35981 ;
  assign n35983 = n35982 ^ n35171 ;
  assign n35979 = n35338 ^ n35337 ;
  assign n35980 = n35979 ^ n35182 ;
  assign n35984 = n35983 ^ n35980 ;
  assign n35985 = ~n34592 & n35984 ;
  assign n35986 = n35985 ^ n35182 ;
  assign n35987 = n35986 ^ n33688 ;
  assign n35991 = n35990 ^ n35987 ;
  assign n35992 = n35991 ^ x58 ;
  assign n35976 = n35972 ^ n35958 ;
  assign n35977 = ~n35973 & n35976 ;
  assign n35978 = n35977 ^ x59 ;
  assign n35993 = n35992 ^ n35978 ;
  assign n35975 = n35955 & ~n35974 ;
  assign n35994 = n35993 ^ n35975 ;
  assign n35995 = n35994 ^ n35538 ;
  assign n36162 = n36087 ^ n35995 ;
  assign n36163 = ~n34982 & ~n36162 ;
  assign n36164 = n36163 ^ n35538 ;
  assign n36371 = n36370 ^ n36164 ;
  assign n36469 = n36371 ^ x278 ;
  assign n36470 = n36469 ^ n36371 ;
  assign n36471 = n36470 ^ n36373 ;
  assign n36472 = ~n36468 & n36471 ;
  assign n36473 = n36472 ^ n36469 ;
  assign n36561 = n36473 ^ x277 ;
  assign n36562 = n36560 & ~n36561 ;
  assign n36372 = n36371 ^ x277 ;
  assign n36474 = ~n36372 & n36473 ;
  assign n36475 = n36474 ^ x277 ;
  assign n36563 = n36475 ^ x276 ;
  assign n36165 = n36164 ^ n34403 ;
  assign n36299 = n36298 ^ n36164 ;
  assign n36300 = ~n36165 & n36299 ;
  assign n36301 = n36300 ^ n34403 ;
  assign n36367 = n36301 ^ n34485 ;
  assign n36112 = n35975 & n35993 ;
  assign n36108 = n35991 ^ n35978 ;
  assign n36109 = n35992 & ~n36108 ;
  assign n36110 = n36109 ^ x58 ;
  assign n36095 = n35983 ^ n35979 ;
  assign n36096 = n35340 ^ n35339 ;
  assign n36097 = n36096 ^ n35182 ;
  assign n36098 = n36097 ^ n35979 ;
  assign n36099 = n36098 ^ n36096 ;
  assign n36100 = ~n36095 & n36099 ;
  assign n36101 = n36100 ^ n36097 ;
  assign n36102 = n36101 ^ n35375 ;
  assign n36103 = n34712 & ~n36102 ;
  assign n36104 = n36103 ^ n35375 ;
  assign n36105 = n36104 ^ n33887 ;
  assign n36091 = n35990 ^ n35986 ;
  assign n36092 = n35990 ^ n33688 ;
  assign n36093 = ~n36091 & n36092 ;
  assign n36094 = n36093 ^ n33688 ;
  assign n36106 = n36105 ^ n36094 ;
  assign n36107 = n36106 ^ x57 ;
  assign n36111 = n36110 ^ n36107 ;
  assign n36113 = n36112 ^ n36111 ;
  assign n36302 = n36113 ^ n35534 ;
  assign n36088 = n36087 ^ n35994 ;
  assign n36089 = n35995 & ~n36088 ;
  assign n36090 = n36089 ^ n35538 ;
  assign n36303 = n36302 ^ n36090 ;
  assign n36304 = ~n35124 & n36303 ;
  assign n36305 = n36304 ^ n35534 ;
  assign n36368 = n36367 ^ n36305 ;
  assign n36564 = n36563 ^ n36368 ;
  assign n36565 = ~n36562 & n36564 ;
  assign n36369 = n36368 ^ x276 ;
  assign n36476 = n36475 ^ n36368 ;
  assign n36477 = ~n36369 & n36476 ;
  assign n36478 = n36477 ^ x276 ;
  assign n36306 = n36305 ^ n36301 ;
  assign n36310 = ~n36306 & ~n36367 ;
  assign n36114 = n36113 ^ n36090 ;
  assign n36132 = n36104 ^ n36094 ;
  assign n36133 = n36105 & n36132 ;
  assign n36129 = n35467 ^ n33887 ;
  assign n36130 = n36129 ^ n33903 ;
  assign n36131 = n36130 ^ x56 ;
  assign n36134 = n36133 ^ n36131 ;
  assign n36125 = n36096 ^ n35375 ;
  assign n36126 = n36101 & ~n36125 ;
  assign n36122 = n35342 ^ n35341 ;
  assign n36123 = n36122 ^ n35467 ;
  assign n36124 = n36123 ^ n36096 ;
  assign n36127 = n36126 ^ n36124 ;
  assign n36128 = ~n34778 & n36127 ;
  assign n36135 = n36134 ^ n36128 ;
  assign n36115 = n36112 ^ n36110 ;
  assign n36117 = n36110 ^ n36106 ;
  assign n36120 = ~n36115 & ~n36117 ;
  assign n36118 = n36117 ^ n36112 ;
  assign n36119 = ~x57 & n36118 ;
  assign n36121 = n36120 ^ n36119 ;
  assign n36136 = n36135 ^ n36121 ;
  assign n36137 = n36136 ^ n35534 ;
  assign n36138 = n36137 ^ n36090 ;
  assign n36139 = n36138 ^ n36136 ;
  assign n36140 = ~n36114 & ~n36139 ;
  assign n36141 = n36140 ^ n36137 ;
  assign n36158 = n36141 ^ n35677 ;
  assign n36159 = n34978 & ~n36158 ;
  assign n36160 = n36159 ^ n35677 ;
  assign n36307 = n36160 ^ n34485 ;
  assign n36311 = n36310 ^ n36307 ;
  assign n36365 = n36311 ^ n34543 ;
  assign n36366 = n36365 ^ x275 ;
  assign n36566 = n36478 ^ n36366 ;
  assign n36567 = ~n36565 & ~n36566 ;
  assign n36479 = n36478 ^ n36365 ;
  assign n36480 = ~n36366 & n36479 ;
  assign n36481 = n36480 ^ x275 ;
  assign n36161 = n36160 ^ n34543 ;
  assign n36312 = n36161 & ~n36311 ;
  assign n36313 = n36312 ^ n34543 ;
  assign n36362 = n36313 ^ n34401 ;
  assign n36144 = n35677 ^ n35512 ;
  assign n36142 = n36136 ^ n35677 ;
  assign n36143 = ~n36141 & ~n36142 ;
  assign n36145 = n36144 ^ n36143 ;
  assign n36154 = n36145 ^ n35508 ;
  assign n36155 = n34975 & ~n36154 ;
  assign n36156 = n36155 ^ n35508 ;
  assign n36363 = n36362 ^ n36156 ;
  assign n36364 = n36363 ^ x274 ;
  assign n36568 = n36481 ^ n36364 ;
  assign n36569 = ~n36567 & n36568 ;
  assign n36482 = n36481 ^ n36363 ;
  assign n36483 = ~n36364 & n36482 ;
  assign n36484 = n36483 ^ x274 ;
  assign n36570 = n36484 ^ x273 ;
  assign n36157 = n36156 ^ n34401 ;
  assign n36314 = n36313 ^ n36156 ;
  assign n36315 = n36157 & n36314 ;
  assign n36316 = n36315 ^ n34401 ;
  assign n36148 = n35852 ^ n35512 ;
  assign n36149 = n36148 ^ n35529 ;
  assign n35513 = n35512 ^ n35508 ;
  assign n36146 = n35513 & ~n36145 ;
  assign n36147 = n36146 ^ n35512 ;
  assign n36150 = n36149 ^ n36147 ;
  assign n36151 = n34884 & n36150 ;
  assign n36152 = n36151 ^ n35529 ;
  assign n36153 = n36152 ^ n34478 ;
  assign n36360 = n36316 ^ n36153 ;
  assign n36571 = n36570 ^ n36360 ;
  assign n36572 = ~n36569 & ~n36571 ;
  assign n36361 = n36360 ^ x273 ;
  assign n36485 = n36484 ^ n36360 ;
  assign n36486 = ~n36361 & n36485 ;
  assign n36487 = n36486 ^ x273 ;
  assign n36317 = n36316 ^ n36152 ;
  assign n36318 = ~n36153 & ~n36317 ;
  assign n36319 = n36318 ^ n34478 ;
  assign n36357 = n36319 ^ n34474 ;
  assign n36323 = n35854 ^ n35853 ;
  assign n36324 = n36323 ^ n35526 ;
  assign n36320 = n36147 ^ n35529 ;
  assign n36321 = n36149 & ~n36320 ;
  assign n36322 = n36321 ^ n36148 ;
  assign n36325 = n36324 ^ n36322 ;
  assign n36326 = n35026 & ~n36325 ;
  assign n36327 = n36326 ^ n35526 ;
  assign n36358 = n36357 ^ n36327 ;
  assign n36359 = n36358 ^ x272 ;
  assign n36573 = n36487 ^ n36359 ;
  assign n36574 = ~n36572 & n36573 ;
  assign n36488 = n36487 ^ n36358 ;
  assign n36489 = ~n36359 & n36488 ;
  assign n36490 = n36489 ^ x272 ;
  assign n36575 = n36490 ^ x287 ;
  assign n36328 = n36327 ^ n36319 ;
  assign n36332 = n35857 ^ n35855 ;
  assign n36333 = n36332 ^ n35827 ;
  assign n36329 = n36322 ^ n35526 ;
  assign n36330 = ~n36324 & ~n36329 ;
  assign n36331 = n36330 ^ n36323 ;
  assign n36334 = n36333 ^ n36331 ;
  assign n36335 = ~n35147 & ~n36334 ;
  assign n36336 = n36335 ^ n35827 ;
  assign n36337 = n36336 ^ n34474 ;
  assign n36338 = n36337 ^ n36319 ;
  assign n36339 = n36338 ^ n36336 ;
  assign n36340 = n36328 & ~n36339 ;
  assign n36341 = n36340 ^ n36337 ;
  assign n36491 = n36341 ^ n34560 ;
  assign n36576 = n36575 ^ n36491 ;
  assign n36577 = n36574 & n36576 ;
  assign n36492 = n36491 ^ n36490 ;
  assign n36345 = n35859 ^ n35858 ;
  assign n36346 = n36345 ^ n35905 ;
  assign n36342 = n36331 ^ n35827 ;
  assign n36343 = n36333 & n36342 ;
  assign n36344 = n36343 ^ n36332 ;
  assign n36347 = n36346 ^ n36344 ;
  assign n36348 = n35022 & n36347 ;
  assign n36349 = n36348 ^ n35905 ;
  assign n36351 = n36349 ^ n34560 ;
  assign n36350 = n36349 ^ n36336 ;
  assign n36352 = n36351 ^ n36350 ;
  assign n36353 = ~n36341 & ~n36352 ;
  assign n36354 = n36353 ^ n36351 ;
  assign n36355 = n36354 ^ n34470 ;
  assign n36493 = n36355 ^ x287 ;
  assign n36494 = n36493 ^ n36355 ;
  assign n36495 = n36494 ^ n36490 ;
  assign n36496 = n36492 & n36495 ;
  assign n36497 = n36496 ^ n36493 ;
  assign n36578 = n36497 ^ x286 ;
  assign n36579 = n36577 & n36578 ;
  assign n36508 = n35861 ^ n35860 ;
  assign n36506 = n36345 ^ n35929 ;
  assign n36504 = n36344 ^ n35905 ;
  assign n36505 = n36346 & n36504 ;
  assign n36507 = n36506 ^ n36505 ;
  assign n36509 = n36508 ^ n36507 ;
  assign n36510 = n35018 & n36509 ;
  assign n36511 = n36510 ^ n35929 ;
  assign n36512 = n36511 ^ n34466 ;
  assign n36501 = n36349 ^ n34470 ;
  assign n36502 = ~n36354 & n36501 ;
  assign n36503 = n36502 ^ n34470 ;
  assign n36513 = n36512 ^ n36503 ;
  assign n36356 = n36355 ^ x286 ;
  assign n36498 = ~n36356 & n36497 ;
  assign n36499 = n36498 ^ x286 ;
  assign n36500 = n36499 ^ x285 ;
  assign n36514 = n36513 ^ n36500 ;
  assign n36580 = n36579 ^ n36514 ;
  assign n36581 = n36580 ^ n36209 ;
  assign n37684 = n36580 ^ n36015 ;
  assign n36793 = n36547 ^ n36545 ;
  assign n36788 = n36303 ^ n36162 ;
  assign n36740 = n36542 ^ n36540 ;
  assign n36741 = n36740 ^ n36167 ;
  assign n36743 = n36536 ^ n36535 ;
  assign n36744 = n36743 ^ n36171 ;
  assign n36745 = n36534 ^ n36532 ;
  assign n36746 = n36745 ^ n36175 ;
  assign n36747 = n36531 ^ n36515 ;
  assign n36748 = n36747 ^ n36179 ;
  assign n36750 = n36527 ^ n36526 ;
  assign n36751 = n36750 ^ n36182 ;
  assign n36752 = n36525 ^ n36516 ;
  assign n36753 = n36752 ^ n36186 ;
  assign n36732 = n36524 ^ n36523 ;
  assign n36756 = n36732 ^ n36186 ;
  assign n36733 = n36732 ^ n36190 ;
  assign n36582 = n36522 ^ n36520 ;
  assign n36583 = n36582 ^ n36195 ;
  assign n36584 = n36519 ^ n36517 ;
  assign n36585 = n36584 ^ n36198 ;
  assign n36586 = n36508 ^ n35929 ;
  assign n36587 = ~n36507 & ~n36586 ;
  assign n36588 = n36587 ^ n36508 ;
  assign n36602 = n36588 ^ n35948 ;
  assign n36603 = n35865 ^ n35864 ;
  assign n36589 = n35863 ^ n35862 ;
  assign n36604 = n36603 ^ n36589 ;
  assign n36605 = n36604 ^ n36603 ;
  assign n36606 = n36605 ^ n36588 ;
  assign n36607 = ~n36602 & ~n36606 ;
  assign n36608 = n36607 ^ n36604 ;
  assign n36609 = n36608 ^ n35965 ;
  assign n36610 = ~n35171 & ~n36609 ;
  assign n36611 = n36610 ^ n35965 ;
  assign n36590 = n36589 ^ n35948 ;
  assign n36591 = n36590 ^ n36588 ;
  assign n36592 = ~n35014 & ~n36591 ;
  assign n36593 = n36592 ^ n35948 ;
  assign n36594 = n36593 ^ n34575 ;
  assign n36595 = n36511 ^ n36503 ;
  assign n36596 = n36512 & ~n36595 ;
  assign n36597 = n36596 ^ n34466 ;
  assign n36598 = n36597 ^ n36593 ;
  assign n36599 = ~n36594 & n36598 ;
  assign n36600 = n36599 ^ n34575 ;
  assign n36627 = n36611 ^ n36600 ;
  assign n36628 = n35868 ^ n35866 ;
  assign n36630 = n36628 ^ n35965 ;
  assign n36629 = n36628 ^ n36603 ;
  assign n36631 = n36630 ^ n36629 ;
  assign n36632 = ~n36608 & n36631 ;
  assign n36633 = n36632 ^ n36630 ;
  assign n36634 = n36633 ^ n35984 ;
  assign n36635 = ~n35182 & n36634 ;
  assign n36636 = n36635 ^ n35984 ;
  assign n36637 = n36636 ^ n34463 ;
  assign n36638 = n36637 ^ n36600 ;
  assign n36639 = n36638 ^ n36636 ;
  assign n36640 = ~n36627 & n36639 ;
  assign n36641 = n36640 ^ n36637 ;
  assign n36642 = n36641 ^ n34592 ;
  assign n36601 = n36600 ^ n34463 ;
  assign n36612 = n36611 ^ n36601 ;
  assign n36613 = n36612 ^ x283 ;
  assign n36614 = n36597 ^ n34575 ;
  assign n36615 = n36614 ^ n36593 ;
  assign n36616 = n36615 ^ x284 ;
  assign n36617 = n36513 ^ x285 ;
  assign n36618 = n36513 ^ n36499 ;
  assign n36619 = ~n36617 & n36618 ;
  assign n36620 = n36619 ^ x285 ;
  assign n36621 = n36620 ^ n36615 ;
  assign n36622 = n36616 & ~n36621 ;
  assign n36623 = n36622 ^ x284 ;
  assign n36624 = n36623 ^ n36612 ;
  assign n36625 = ~n36613 & n36624 ;
  assign n36626 = n36625 ^ x283 ;
  assign n36643 = n36642 ^ n36626 ;
  assign n36654 = n36636 ^ n34592 ;
  assign n36655 = n36641 & ~n36654 ;
  assign n36656 = n36655 ^ n34592 ;
  assign n36644 = n35870 ^ n35869 ;
  assign n36646 = n36644 ^ n35984 ;
  assign n36645 = n36644 ^ n36628 ;
  assign n36647 = n36646 ^ n36645 ;
  assign n36648 = ~n36633 & ~n36647 ;
  assign n36649 = n36648 ^ n36646 ;
  assign n36650 = n36649 ^ n36102 ;
  assign n36651 = n35375 & n36650 ;
  assign n36652 = n36651 ^ n36102 ;
  assign n36653 = n36652 ^ n34712 ;
  assign n36657 = n36656 ^ n36653 ;
  assign n36658 = n36657 ^ x282 ;
  assign n36659 = n36658 ^ n36626 ;
  assign n36660 = n36659 ^ n36657 ;
  assign n36661 = ~n36643 & n36660 ;
  assign n36662 = n36661 ^ n36658 ;
  assign n36693 = n36662 ^ x281 ;
  assign n36664 = n36514 & n36579 ;
  assign n36665 = n36620 ^ n36616 ;
  assign n36666 = n36664 & ~n36665 ;
  assign n36667 = n36623 ^ n36613 ;
  assign n36668 = ~n36666 & ~n36667 ;
  assign n36669 = n36642 ^ x282 ;
  assign n36670 = n36669 ^ n36626 ;
  assign n36671 = ~n36668 & ~n36670 ;
  assign n36694 = n36693 ^ n36671 ;
  assign n36695 = n36694 ^ n36230 ;
  assign n36702 = n36667 ^ n36666 ;
  assign n36696 = ~n36209 & ~n36580 ;
  assign n36697 = n36696 ^ n36214 ;
  assign n36698 = n36665 ^ n36664 ;
  assign n36699 = n36698 ^ n36696 ;
  assign n36700 = ~n36697 & ~n36699 ;
  assign n36701 = n36700 ^ n36214 ;
  assign n36703 = n36702 ^ n36701 ;
  assign n36704 = n36670 ^ n36668 ;
  assign n36705 = n36704 ^ n36205 ;
  assign n36706 = n36705 ^ n36701 ;
  assign n36707 = n36706 ^ n36704 ;
  assign n36708 = n36703 & ~n36707 ;
  assign n36709 = n36708 ^ n36705 ;
  assign n36711 = n36694 ^ n36203 ;
  assign n36710 = n36704 ^ n36694 ;
  assign n36712 = n36711 ^ n36710 ;
  assign n36713 = n36709 & ~n36712 ;
  assign n36714 = n36713 ^ n36711 ;
  assign n36715 = ~n36695 & ~n36714 ;
  assign n36716 = n36715 ^ n36230 ;
  assign n36687 = n36644 ^ n36102 ;
  assign n36688 = ~n36649 & n36687 ;
  assign n36684 = n35872 ^ n35871 ;
  assign n36685 = n36684 ^ n36127 ;
  assign n36686 = n36685 ^ n36644 ;
  assign n36689 = n36688 ^ n36686 ;
  assign n36690 = n35467 & n36689 ;
  assign n36680 = n34778 ^ n34712 ;
  assign n36681 = n36680 ^ n36127 ;
  assign n36682 = n36681 ^ x280 ;
  assign n36677 = n36656 ^ n36652 ;
  assign n36678 = n36656 ^ n34712 ;
  assign n36679 = ~n36677 & ~n36678 ;
  assign n36683 = n36682 ^ n36679 ;
  assign n36691 = n36690 ^ n36683 ;
  assign n36672 = n36671 ^ n36657 ;
  assign n36675 = ~n36662 & n36672 ;
  assign n36663 = n36662 ^ n36657 ;
  assign n36673 = n36672 ^ n36663 ;
  assign n36674 = x281 & n36673 ;
  assign n36676 = n36675 ^ n36674 ;
  assign n36692 = n36691 ^ n36676 ;
  assign n36717 = n36716 ^ n36692 ;
  assign n36718 = n36716 ^ n36237 ;
  assign n36719 = n36717 & ~n36718 ;
  assign n36720 = n36719 ^ n36237 ;
  assign n36721 = n36720 ^ n36245 ;
  assign n36724 = n36720 ^ n36517 ;
  assign n36725 = ~n36721 & ~n36724 ;
  assign n36722 = n36517 ^ n36198 ;
  assign n36726 = n36725 ^ n36722 ;
  assign n36727 = n36585 & ~n36726 ;
  assign n36728 = n36727 ^ n36584 ;
  assign n36729 = n36728 ^ n36195 ;
  assign n36730 = ~n36583 & n36729 ;
  assign n36731 = n36730 ^ n36582 ;
  assign n36754 = n36731 ^ n36190 ;
  assign n36755 = n36733 & ~n36754 ;
  assign n36757 = n36756 ^ n36755 ;
  assign n36758 = ~n36753 & n36757 ;
  assign n36759 = n36758 ^ n36752 ;
  assign n36760 = n36759 ^ n36750 ;
  assign n36761 = ~n36751 & n36760 ;
  assign n36762 = n36761 ^ n36182 ;
  assign n36749 = n36530 ^ n36528 ;
  assign n36763 = n36762 ^ n36749 ;
  assign n36764 = n36747 ^ n36271 ;
  assign n36765 = n36764 ^ n36749 ;
  assign n36766 = n36765 ^ n36747 ;
  assign n36767 = ~n36763 & n36766 ;
  assign n36768 = n36767 ^ n36764 ;
  assign n36769 = n36748 & ~n36768 ;
  assign n36770 = n36769 ^ n36179 ;
  assign n36771 = n36770 ^ n36745 ;
  assign n36772 = ~n36746 & ~n36771 ;
  assign n36773 = n36772 ^ n36175 ;
  assign n36774 = n36773 ^ n36743 ;
  assign n36775 = n36744 & ~n36774 ;
  assign n36776 = n36775 ^ n36171 ;
  assign n36742 = n36539 ^ n36537 ;
  assign n36777 = n36776 ^ n36742 ;
  assign n36779 = n36740 ^ n36288 ;
  assign n36778 = n36776 ^ n36740 ;
  assign n36780 = n36779 ^ n36778 ;
  assign n36781 = ~n36777 & n36780 ;
  assign n36782 = n36781 ^ n36779 ;
  assign n36783 = n36741 & ~n36782 ;
  assign n36739 = n36167 ^ n36162 ;
  assign n36784 = n36783 ^ n36739 ;
  assign n36785 = n36544 ^ n36543 ;
  assign n36786 = n36785 ^ n36162 ;
  assign n36787 = n36784 & ~n36786 ;
  assign n36789 = n36788 ^ n36787 ;
  assign n36989 = n36793 ^ n36789 ;
  assign n37082 = ~n35534 & n36989 ;
  assign n37083 = n37082 ^ n36303 ;
  assign n37084 = n37083 ^ n35124 ;
  assign n36992 = n36785 ^ n36784 ;
  assign n37121 = n35538 & n36992 ;
  assign n37122 = n37121 ^ n36162 ;
  assign n36996 = n36782 ^ n36167 ;
  assign n37085 = n35542 & ~n36996 ;
  assign n37086 = n37085 ^ n36167 ;
  assign n37087 = n37086 ^ n34985 ;
  assign n36998 = n36777 ^ n36288 ;
  assign n37088 = ~n35547 & ~n36998 ;
  assign n37089 = n37088 ^ n36288 ;
  assign n37090 = n37089 ^ n35107 ;
  assign n37001 = n36773 ^ n36744 ;
  assign n37091 = n35551 & ~n37001 ;
  assign n37092 = n37091 ^ n36171 ;
  assign n37093 = n37092 ^ n35038 ;
  assign n37009 = n36768 ^ n36179 ;
  assign n37098 = ~n35555 & n37009 ;
  assign n37099 = n37098 ^ n36179 ;
  assign n36886 = n36759 ^ n36751 ;
  assign n36887 = ~n35563 & ~n36886 ;
  assign n36888 = n36887 ^ n36182 ;
  assign n36959 = n36888 ^ n35080 ;
  assign n36805 = n36757 ^ n36752 ;
  assign n36806 = n35636 & ~n36805 ;
  assign n36807 = n36806 ^ n36186 ;
  assign n36808 = n36807 ^ n35047 ;
  assign n36734 = n36733 ^ n36731 ;
  assign n36809 = n35629 & n36734 ;
  assign n36810 = n36809 ^ n36190 ;
  assign n36811 = n36810 ^ n35051 ;
  assign n36815 = n36517 ^ n36245 ;
  assign n36816 = n36815 ^ n36720 ;
  assign n36817 = ~n35576 & n36816 ;
  assign n36818 = n36817 ^ n36245 ;
  assign n36819 = n36818 ^ n34885 ;
  assign n36854 = n36692 ^ n36237 ;
  assign n36855 = n36854 ^ n36716 ;
  assign n36856 = n35581 & n36855 ;
  assign n36857 = n36856 ^ n36237 ;
  assign n36820 = n36714 ^ n36230 ;
  assign n36821 = n35609 & n36820 ;
  assign n36822 = n36821 ^ n36230 ;
  assign n36823 = n36822 ^ n34892 ;
  assign n36828 = n35509 & ~n36581 ;
  assign n36829 = n36828 ^ n36209 ;
  assign n36830 = ~n34904 & n36829 ;
  assign n36831 = n36830 ^ n34909 ;
  assign n36832 = n36698 ^ n36697 ;
  assign n36833 = ~n35591 & n36832 ;
  assign n36834 = n36833 ^ n36214 ;
  assign n36835 = n36834 ^ n36830 ;
  assign n36836 = n36831 & ~n36835 ;
  assign n36837 = n36836 ^ n34909 ;
  assign n36824 = n36701 ^ n36205 ;
  assign n36825 = n36824 ^ n36702 ;
  assign n36826 = n35600 & n36825 ;
  assign n36827 = n36826 ^ n36205 ;
  assign n36838 = n36837 ^ n36827 ;
  assign n36839 = n36709 ^ n36203 ;
  assign n36840 = n35585 & n36839 ;
  assign n36841 = n36840 ^ n36203 ;
  assign n36842 = n36841 ^ n34900 ;
  assign n36843 = n36842 ^ n36827 ;
  assign n36844 = n36843 ^ n36841 ;
  assign n36845 = n36838 & n36844 ;
  assign n36846 = n36845 ^ n36842 ;
  assign n36848 = n36822 ^ n34896 ;
  assign n36847 = n36841 ^ n36822 ;
  assign n36849 = n36848 ^ n36847 ;
  assign n36850 = ~n36846 & n36849 ;
  assign n36851 = n36850 ^ n36848 ;
  assign n36852 = ~n36823 & n36851 ;
  assign n36853 = n36852 ^ n34892 ;
  assign n36858 = n36857 ^ n36853 ;
  assign n36859 = n36818 ^ n34888 ;
  assign n36860 = n36859 ^ n36818 ;
  assign n36861 = n36860 ^ n36853 ;
  assign n36862 = ~n36858 & n36861 ;
  assign n36863 = n36862 ^ n36859 ;
  assign n36864 = n36819 & ~n36863 ;
  assign n36865 = n36864 ^ n34885 ;
  assign n36812 = n36726 ^ n36584 ;
  assign n36813 = ~n35571 & n36812 ;
  assign n36814 = n36813 ^ n36198 ;
  assign n36866 = n36865 ^ n36814 ;
  assign n36867 = n36728 ^ n36583 ;
  assign n36868 = ~n35566 & ~n36867 ;
  assign n36869 = n36868 ^ n36195 ;
  assign n36870 = n36869 ^ n35055 ;
  assign n36871 = n36870 ^ n36814 ;
  assign n36872 = n36871 ^ n36869 ;
  assign n36873 = n36866 & ~n36872 ;
  assign n36874 = n36873 ^ n36870 ;
  assign n36876 = n36810 ^ n35065 ;
  assign n36875 = n36869 ^ n36810 ;
  assign n36877 = n36876 ^ n36875 ;
  assign n36878 = ~n36874 & n36877 ;
  assign n36879 = n36878 ^ n36876 ;
  assign n36880 = ~n36811 & n36879 ;
  assign n36881 = n36880 ^ n35051 ;
  assign n36882 = n36881 ^ n36807 ;
  assign n36883 = ~n36808 & ~n36882 ;
  assign n36884 = n36883 ^ n35047 ;
  assign n36960 = n36888 ^ n36884 ;
  assign n36961 = n36959 & ~n36960 ;
  assign n36962 = n36961 ^ n35080 ;
  assign n36954 = n36749 ^ n36271 ;
  assign n36955 = n36954 ^ n36762 ;
  assign n36956 = ~n35559 & n36955 ;
  assign n36957 = n36956 ^ n36271 ;
  assign n37094 = n36962 ^ n36957 ;
  assign n37095 = n36962 ^ n35043 ;
  assign n37096 = ~n37094 & ~n37095 ;
  assign n37097 = n37096 ^ n35043 ;
  assign n37100 = n37099 ^ n37097 ;
  assign n37003 = n36770 ^ n36746 ;
  assign n37101 = n35653 & ~n37003 ;
  assign n37102 = n37101 ^ n36175 ;
  assign n37103 = n37102 ^ n35091 ;
  assign n37104 = n37103 ^ n37102 ;
  assign n37105 = n37104 ^ n37097 ;
  assign n37106 = n37100 & n37105 ;
  assign n37107 = n37106 ^ n37103 ;
  assign n37109 = n37092 ^ n35097 ;
  assign n37108 = n37102 ^ n37092 ;
  assign n37110 = n37109 ^ n37108 ;
  assign n37111 = ~n37107 & n37110 ;
  assign n37112 = n37111 ^ n37109 ;
  assign n37113 = ~n37093 & ~n37112 ;
  assign n37114 = n37113 ^ n35038 ;
  assign n37115 = n37114 ^ n37089 ;
  assign n37116 = n37090 & n37115 ;
  assign n37117 = n37116 ^ n35107 ;
  assign n37118 = n37117 ^ n37086 ;
  assign n37119 = ~n37087 & ~n37118 ;
  assign n37120 = n37119 ^ n34985 ;
  assign n37123 = n37122 ^ n37120 ;
  assign n37124 = n37083 ^ n34982 ;
  assign n37125 = n37124 ^ n37083 ;
  assign n37126 = n37125 ^ n37120 ;
  assign n37127 = n37123 & ~n37126 ;
  assign n37128 = n37127 ^ n37124 ;
  assign n37129 = ~n37084 & n37128 ;
  assign n37130 = n37129 ^ n35124 ;
  assign n37178 = n37130 ^ n34978 ;
  assign n36790 = n36550 ^ n36548 ;
  assign n36791 = n36790 ^ n36303 ;
  assign n36792 = n36791 ^ n36790 ;
  assign n36794 = n36793 ^ n36792 ;
  assign n36795 = ~n36789 & ~n36794 ;
  assign n36796 = n36795 ^ n36791 ;
  assign n36986 = n36796 ^ n36158 ;
  assign n37079 = n35677 & n36986 ;
  assign n37080 = n37079 ^ n36158 ;
  assign n37179 = n37178 ^ n37080 ;
  assign n37180 = n37179 ^ x499 ;
  assign n37181 = n37120 ^ n34982 ;
  assign n37182 = n37181 ^ n37122 ;
  assign n37183 = n37182 ^ x501 ;
  assign n37184 = n37117 ^ n34985 ;
  assign n37185 = n37184 ^ n37086 ;
  assign n37186 = n37185 ^ x502 ;
  assign n37207 = n37114 ^ n37090 ;
  assign n37187 = n37112 ^ n35038 ;
  assign n37188 = n37187 ^ x488 ;
  assign n37189 = n37107 ^ n35097 ;
  assign n37190 = n37189 ^ x489 ;
  assign n36958 = n36957 ^ n35043 ;
  assign n36963 = n36962 ^ n36958 ;
  assign n37193 = n36963 ^ x491 ;
  assign n36885 = n36884 ^ n35080 ;
  assign n36889 = n36888 ^ n36885 ;
  assign n36890 = n36889 ^ x492 ;
  assign n36891 = n36881 ^ n36808 ;
  assign n36892 = n36891 ^ x493 ;
  assign n36894 = n36814 ^ n35055 ;
  assign n36895 = n36894 ^ n36865 ;
  assign n36896 = n36895 ^ x480 ;
  assign n36898 = n36857 ^ n34888 ;
  assign n36899 = n36898 ^ n36853 ;
  assign n36900 = n36899 ^ x482 ;
  assign n36901 = n36851 ^ n34892 ;
  assign n36902 = n36901 ^ x483 ;
  assign n36904 = n36837 ^ n34900 ;
  assign n36905 = n36904 ^ n36827 ;
  assign n36906 = n36905 ^ x485 ;
  assign n36908 = n36015 ^ n35395 ;
  assign n36909 = n36908 ^ n36828 ;
  assign n36910 = x487 & ~n36909 ;
  assign n36907 = n36834 ^ n36831 ;
  assign n36911 = n36910 ^ n36907 ;
  assign n36912 = n36905 ^ x486 ;
  assign n36913 = n36912 ^ n36905 ;
  assign n36914 = n36913 ^ n36907 ;
  assign n36915 = ~n36911 & n36914 ;
  assign n36916 = n36915 ^ n36912 ;
  assign n36917 = n36906 & ~n36916 ;
  assign n36918 = n36917 ^ x485 ;
  assign n36903 = n36846 ^ n34896 ;
  assign n36919 = n36918 ^ n36903 ;
  assign n36920 = n36918 ^ x484 ;
  assign n36921 = n36919 & n36920 ;
  assign n36922 = n36921 ^ x484 ;
  assign n36923 = n36922 ^ n36901 ;
  assign n36924 = n36902 & ~n36923 ;
  assign n36925 = n36924 ^ x483 ;
  assign n36926 = n36925 ^ n36899 ;
  assign n36927 = ~n36900 & n36926 ;
  assign n36928 = n36927 ^ x482 ;
  assign n36897 = n36863 ^ n34885 ;
  assign n36929 = n36928 ^ n36897 ;
  assign n36930 = n36928 ^ x481 ;
  assign n36931 = n36929 & n36930 ;
  assign n36932 = n36931 ^ x481 ;
  assign n36933 = n36932 ^ n36895 ;
  assign n36934 = n36896 & ~n36933 ;
  assign n36935 = n36934 ^ x480 ;
  assign n36893 = n36874 ^ n35065 ;
  assign n36936 = n36935 ^ n36893 ;
  assign n36937 = n36879 ^ n35051 ;
  assign n36938 = n36937 ^ x495 ;
  assign n36939 = n36938 ^ n36893 ;
  assign n36940 = n36939 ^ n36937 ;
  assign n36941 = n36936 & ~n36940 ;
  assign n36942 = n36941 ^ n36938 ;
  assign n36944 = n36891 ^ x494 ;
  assign n36943 = n36937 ^ n36891 ;
  assign n36945 = n36944 ^ n36943 ;
  assign n36946 = ~n36942 & n36945 ;
  assign n36947 = n36946 ^ n36944 ;
  assign n36948 = n36892 & ~n36947 ;
  assign n36949 = n36948 ^ x493 ;
  assign n36950 = n36949 ^ n36889 ;
  assign n36951 = n36890 & ~n36950 ;
  assign n36952 = n36951 ^ x492 ;
  assign n37194 = n36963 ^ n36952 ;
  assign n37195 = ~n37193 & n37194 ;
  assign n37196 = n37195 ^ x491 ;
  assign n37191 = n37099 ^ n35091 ;
  assign n37192 = n37191 ^ n37097 ;
  assign n37197 = n37196 ^ n37192 ;
  assign n37198 = n37196 ^ x490 ;
  assign n37199 = ~n37197 & n37198 ;
  assign n37200 = n37199 ^ x490 ;
  assign n37201 = n37200 ^ n37189 ;
  assign n37202 = ~n37190 & n37201 ;
  assign n37203 = n37202 ^ x489 ;
  assign n37204 = n37203 ^ n37187 ;
  assign n37205 = n37188 & ~n37204 ;
  assign n37206 = n37205 ^ x488 ;
  assign n37208 = n37207 ^ n37206 ;
  assign n37209 = n37185 ^ x503 ;
  assign n37210 = n37209 ^ n37185 ;
  assign n37211 = n37210 ^ n37206 ;
  assign n37212 = ~n37208 & n37211 ;
  assign n37213 = n37212 ^ n37209 ;
  assign n37214 = n37186 & ~n37213 ;
  assign n37215 = n37214 ^ x502 ;
  assign n37216 = n37215 ^ n37182 ;
  assign n37217 = n37183 & ~n37216 ;
  assign n37218 = n37217 ^ x501 ;
  assign n37219 = n37218 ^ x500 ;
  assign n37220 = n37128 ^ n35124 ;
  assign n37221 = n37220 ^ n37218 ;
  assign n37222 = n37219 & ~n37221 ;
  assign n37223 = n37222 ^ x500 ;
  assign n37224 = n37223 ^ n37179 ;
  assign n37225 = n37180 & ~n37224 ;
  assign n37226 = n37225 ^ x499 ;
  assign n36737 = n36553 ^ n36551 ;
  assign n36798 = n36737 ^ n36158 ;
  assign n36797 = n36790 ^ n36737 ;
  assign n36799 = n36798 ^ n36797 ;
  assign n36800 = n36796 & n36799 ;
  assign n36801 = n36800 ^ n36798 ;
  assign n36983 = n36801 ^ n36154 ;
  assign n37134 = ~n35508 & n36983 ;
  assign n37135 = n37134 ^ n36154 ;
  assign n37176 = n37135 ^ n34975 ;
  assign n37081 = n37080 ^ n34978 ;
  assign n37131 = n37130 ^ n37080 ;
  assign n37132 = ~n37081 & ~n37131 ;
  assign n37133 = n37132 ^ n34978 ;
  assign n37177 = n37176 ^ n37133 ;
  assign n37227 = n37226 ^ n37177 ;
  assign n37136 = n37135 ^ n37133 ;
  assign n36738 = n36737 ^ n36154 ;
  assign n36802 = ~n36738 & n36801 ;
  assign n36803 = n36802 ^ n36154 ;
  assign n36735 = n36556 ^ n36554 ;
  assign n36736 = n36735 ^ n36150 ;
  assign n36804 = n36803 ^ n36736 ;
  assign n37076 = ~n35529 & ~n36804 ;
  assign n37077 = n37076 ^ n36150 ;
  assign n37137 = n37077 ^ n34975 ;
  assign n37138 = n37137 ^ n37077 ;
  assign n37139 = n37138 ^ n37133 ;
  assign n37140 = n37136 & n37139 ;
  assign n37141 = n37140 ^ n37137 ;
  assign n37228 = n37141 ^ n34884 ;
  assign n37229 = n37228 ^ x498 ;
  assign n37230 = n37229 ^ n37177 ;
  assign n37231 = n37230 ^ n37228 ;
  assign n37232 = n37227 & ~n37231 ;
  assign n37233 = n37232 ^ n37229 ;
  assign n37310 = n37233 ^ x497 ;
  assign n37286 = n37215 ^ n37183 ;
  assign n37287 = n37192 ^ x490 ;
  assign n37288 = n37287 ^ n37196 ;
  assign n36953 = n36952 ^ x491 ;
  assign n36964 = n36963 ^ n36953 ;
  assign n36965 = n36925 ^ n36900 ;
  assign n36966 = n36897 ^ x481 ;
  assign n36967 = n36966 ^ n36928 ;
  assign n36968 = n36965 & n36967 ;
  assign n36969 = n36932 ^ n36896 ;
  assign n36970 = n36968 & ~n36969 ;
  assign n36971 = n36893 ^ x495 ;
  assign n36972 = n36971 ^ n36935 ;
  assign n36973 = ~n36970 & ~n36972 ;
  assign n36974 = n36942 ^ x494 ;
  assign n36975 = ~n36973 & ~n36974 ;
  assign n36976 = n36947 ^ x493 ;
  assign n36977 = n36975 & ~n36976 ;
  assign n36978 = n36949 ^ x492 ;
  assign n36979 = n36978 ^ n36889 ;
  assign n36980 = ~n36977 & n36979 ;
  assign n37289 = ~n36964 & n36980 ;
  assign n37290 = ~n37288 & ~n37289 ;
  assign n37291 = n37200 ^ x489 ;
  assign n37292 = n37291 ^ n37189 ;
  assign n37293 = n37290 & n37292 ;
  assign n37294 = n37203 ^ x488 ;
  assign n37295 = n37294 ^ n37187 ;
  assign n37296 = n37293 & ~n37295 ;
  assign n37297 = n37207 ^ x503 ;
  assign n37298 = n37297 ^ n37206 ;
  assign n37299 = ~n37296 & n37298 ;
  assign n37300 = n37213 ^ x502 ;
  assign n37301 = n37299 & n37300 ;
  assign n37302 = ~n37286 & ~n37301 ;
  assign n37303 = n37220 ^ n37219 ;
  assign n37304 = n37302 & ~n37303 ;
  assign n37305 = n37223 ^ n37180 ;
  assign n37306 = ~n37304 & n37305 ;
  assign n37307 = n37177 ^ x498 ;
  assign n37308 = n37307 ^ n37226 ;
  assign n37309 = ~n37306 & n37308 ;
  assign n37358 = n37310 ^ n37309 ;
  assign n37526 = n37358 ^ n36581 ;
  assign n37527 = ~n36209 & n37526 ;
  assign n37685 = n37684 ^ n37527 ;
  assign n37686 = x199 & ~n37685 ;
  assign n37078 = n37077 ^ n34884 ;
  assign n37142 = n37078 & ~n37141 ;
  assign n37143 = n37142 ^ n34884 ;
  assign n37025 = n36559 ^ n36557 ;
  assign n37023 = n36325 ^ n36150 ;
  assign n37020 = n36803 ^ n36735 ;
  assign n37021 = n36803 ^ n36150 ;
  assign n37022 = n37020 & ~n37021 ;
  assign n37024 = n37023 ^ n37022 ;
  assign n37072 = n37025 ^ n37024 ;
  assign n37073 = ~n35526 & n37072 ;
  assign n37074 = n37073 ^ n36325 ;
  assign n37075 = n37074 ^ n35026 ;
  assign n37174 = n37143 ^ n37075 ;
  assign n37235 = n37174 ^ x497 ;
  assign n37234 = n37228 ^ n37174 ;
  assign n37236 = n37235 ^ n37234 ;
  assign n37237 = ~n37233 & n37236 ;
  assign n37238 = n37237 ^ n37235 ;
  assign n37312 = n37238 ^ x496 ;
  assign n37311 = ~n37309 & n37310 ;
  assign n37361 = n37312 ^ n37311 ;
  assign n37359 = n36581 & ~n37358 ;
  assign n37360 = n37359 ^ n36832 ;
  assign n37531 = n37361 ^ n37360 ;
  assign n37532 = ~n36214 & ~n37531 ;
  assign n37533 = n37532 ^ n36832 ;
  assign n37528 = n37527 ^ n36581 ;
  assign n37529 = n35509 & ~n37528 ;
  assign n37530 = n37529 ^ n35591 ;
  assign n37683 = n37533 ^ n37530 ;
  assign n37687 = n37686 ^ n37683 ;
  assign n37144 = n37143 ^ n37074 ;
  assign n37145 = ~n37075 & n37144 ;
  assign n37146 = n37145 ^ n35026 ;
  assign n37242 = n37146 ^ n35147 ;
  assign n37026 = n37025 ^ n36325 ;
  assign n37027 = ~n37024 & n37026 ;
  assign n37028 = n37027 ^ n36325 ;
  assign n37018 = n36561 ^ n36560 ;
  assign n37019 = n37018 ^ n36334 ;
  assign n37068 = n37028 ^ n37019 ;
  assign n37069 = ~n35827 & n37068 ;
  assign n37070 = n37069 ^ n36334 ;
  assign n37243 = n37242 ^ n37070 ;
  assign n37175 = n37174 ^ x496 ;
  assign n37239 = ~n37175 & n37238 ;
  assign n37240 = n37239 ^ x496 ;
  assign n37241 = n37240 ^ x511 ;
  assign n37314 = n37243 ^ n37241 ;
  assign n37313 = n37311 & ~n37312 ;
  assign n37357 = n37314 ^ n37313 ;
  assign n37522 = n37357 ^ n36825 ;
  assign n37362 = n37361 ^ n37359 ;
  assign n37363 = ~n37360 & n37362 ;
  assign n37364 = n37363 ^ n36832 ;
  assign n37523 = n37522 ^ n37364 ;
  assign n37524 = n36205 & ~n37523 ;
  assign n37525 = n37524 ^ n36825 ;
  assign n37680 = n37525 ^ n35600 ;
  assign n37534 = n37533 ^ n37529 ;
  assign n37535 = ~n37530 & ~n37534 ;
  assign n37536 = n37535 ^ n35591 ;
  assign n37681 = n37680 ^ n37536 ;
  assign n37688 = n37681 ^ x198 ;
  assign n37689 = n37688 ^ n37681 ;
  assign n37690 = n37689 ^ n37683 ;
  assign n37691 = n37687 & ~n37690 ;
  assign n37692 = n37691 ^ n37688 ;
  assign n37791 = n37692 ^ x197 ;
  assign n37682 = n37681 ^ x197 ;
  assign n37693 = ~n37682 & n37692 ;
  assign n37694 = n37693 ^ x197 ;
  assign n37792 = n37694 ^ x196 ;
  assign n37537 = n37536 ^ n37525 ;
  assign n37538 = n37536 ^ n35600 ;
  assign n37539 = n37537 & ~n37538 ;
  assign n37540 = n37539 ^ n35600 ;
  assign n37365 = n37364 ^ n37357 ;
  assign n37366 = n37364 ^ n36825 ;
  assign n37367 = n37365 & n37366 ;
  assign n37368 = n37367 ^ n36825 ;
  assign n37071 = n37070 ^ n35147 ;
  assign n37147 = n37146 ^ n37070 ;
  assign n37148 = n37071 & n37147 ;
  assign n37149 = n37148 ^ n35147 ;
  assign n37172 = n37149 ^ n35022 ;
  assign n37029 = n37028 ^ n37018 ;
  assign n37030 = ~n37019 & n37029 ;
  assign n37031 = n37030 ^ n36334 ;
  assign n37016 = n36564 ^ n36562 ;
  assign n37017 = n37016 ^ n36347 ;
  assign n37064 = n37031 ^ n37017 ;
  assign n37065 = n35905 & n37064 ;
  assign n37066 = n37065 ^ n36347 ;
  assign n37173 = n37172 ^ n37066 ;
  assign n37316 = n37173 ^ x510 ;
  assign n37244 = n37243 ^ n37240 ;
  assign n37245 = n37241 & ~n37244 ;
  assign n37246 = n37245 ^ x511 ;
  assign n37317 = n37316 ^ n37246 ;
  assign n37315 = n37313 & n37314 ;
  assign n37355 = n37317 ^ n37315 ;
  assign n37356 = n37355 ^ n36839 ;
  assign n37518 = n37368 ^ n37356 ;
  assign n37519 = n36203 & ~n37518 ;
  assign n37520 = n37519 ^ n36839 ;
  assign n37521 = n37520 ^ n35585 ;
  assign n37678 = n37540 ^ n37521 ;
  assign n37793 = n37792 ^ n37678 ;
  assign n37794 = ~n37791 & n37793 ;
  assign n37369 = n37368 ^ n37355 ;
  assign n37370 = ~n37356 & n37369 ;
  assign n37371 = n37370 ^ n36839 ;
  assign n37545 = n37371 ^ n36820 ;
  assign n37247 = n37246 ^ n37173 ;
  assign n37067 = n37066 ^ n35022 ;
  assign n37150 = n37149 ^ n37066 ;
  assign n37151 = n37067 & n37150 ;
  assign n37152 = n37151 ^ n35022 ;
  assign n37169 = n37152 ^ n35018 ;
  assign n37032 = n37031 ^ n37016 ;
  assign n37033 = ~n37017 & ~n37032 ;
  assign n37034 = n37033 ^ n36347 ;
  assign n37015 = n36566 ^ n36565 ;
  assign n37035 = n37034 ^ n37015 ;
  assign n37060 = n37035 ^ n36509 ;
  assign n37061 = n35929 & ~n37060 ;
  assign n37062 = n37061 ^ n36509 ;
  assign n37170 = n37169 ^ n37062 ;
  assign n37248 = n37170 ^ x510 ;
  assign n37249 = n37248 ^ n37170 ;
  assign n37250 = n37249 ^ n37173 ;
  assign n37251 = n37247 & ~n37250 ;
  assign n37252 = n37251 ^ n37248 ;
  assign n37319 = n37252 ^ x509 ;
  assign n37318 = ~n37315 & n37317 ;
  assign n37353 = n37319 ^ n37318 ;
  assign n37546 = n37545 ^ n37353 ;
  assign n37547 = ~n36230 & ~n37546 ;
  assign n37548 = n37547 ^ n36820 ;
  assign n37541 = n37540 ^ n37520 ;
  assign n37542 = n37521 & ~n37541 ;
  assign n37543 = n37542 ^ n35585 ;
  assign n37544 = n37543 ^ n35609 ;
  assign n37677 = n37548 ^ n37544 ;
  assign n37795 = n37677 ^ x195 ;
  assign n37679 = n37678 ^ x196 ;
  assign n37695 = n37694 ^ n37678 ;
  assign n37696 = n37679 & ~n37695 ;
  assign n37697 = n37696 ^ x196 ;
  assign n37796 = n37795 ^ n37697 ;
  assign n37797 = ~n37794 & ~n37796 ;
  assign n37698 = n37697 ^ n37677 ;
  assign n37699 = n37697 ^ x195 ;
  assign n37700 = ~n37698 & n37699 ;
  assign n37701 = n37700 ^ x195 ;
  assign n37063 = n37062 ^ n35018 ;
  assign n37153 = n37152 ^ n37062 ;
  assign n37154 = n37063 & ~n37153 ;
  assign n37155 = n37154 ^ n35018 ;
  assign n37256 = n37155 ^ n35014 ;
  assign n37013 = n36568 ^ n36567 ;
  assign n37037 = n37013 ^ n36509 ;
  assign n37036 = n37034 ^ n37013 ;
  assign n37038 = n37037 ^ n37036 ;
  assign n37039 = n37035 & n37038 ;
  assign n37040 = n37039 ^ n37037 ;
  assign n37156 = n37040 ^ n36591 ;
  assign n37157 = ~n35948 & n37156 ;
  assign n37158 = n37157 ^ n36591 ;
  assign n37257 = n37256 ^ n37158 ;
  assign n37171 = n37170 ^ x509 ;
  assign n37253 = n37171 & ~n37252 ;
  assign n37254 = n37253 ^ x509 ;
  assign n37255 = n37254 ^ x508 ;
  assign n37321 = n37257 ^ n37255 ;
  assign n37320 = n37318 & ~n37319 ;
  assign n37375 = n37321 ^ n37320 ;
  assign n37552 = n37375 ^ n36855 ;
  assign n37354 = n37353 ^ n36820 ;
  assign n37372 = n37371 ^ n37353 ;
  assign n37373 = ~n37354 & n37372 ;
  assign n37374 = n37373 ^ n36820 ;
  assign n37553 = n37552 ^ n37374 ;
  assign n37554 = n36237 & ~n37553 ;
  assign n37555 = n37554 ^ n36855 ;
  assign n37674 = n37555 ^ n35581 ;
  assign n37549 = n37548 ^ n37543 ;
  assign n37550 = n37544 & ~n37549 ;
  assign n37551 = n37550 ^ n35609 ;
  assign n37675 = n37674 ^ n37551 ;
  assign n37676 = n37675 ^ x194 ;
  assign n37798 = n37701 ^ n37676 ;
  assign n37799 = ~n37797 & n37798 ;
  assign n37556 = n37555 ^ n37551 ;
  assign n37376 = n37375 ^ n37374 ;
  assign n37159 = n37158 ^ n37155 ;
  assign n37043 = n36571 ^ n36569 ;
  assign n37055 = n37043 ^ n36609 ;
  assign n37014 = n37013 ^ n36591 ;
  assign n37041 = n37014 & n37040 ;
  assign n37042 = n37041 ^ n36591 ;
  assign n37056 = n37055 ^ n37042 ;
  assign n37057 = n35965 & ~n37056 ;
  assign n37058 = n37057 ^ n36609 ;
  assign n37160 = n37058 ^ n35014 ;
  assign n37161 = n37160 ^ n37058 ;
  assign n37162 = n37161 ^ n37155 ;
  assign n37163 = n37159 & ~n37162 ;
  assign n37164 = n37163 ^ n37160 ;
  assign n37262 = n37164 ^ n35171 ;
  assign n37258 = n37257 ^ n37254 ;
  assign n37259 = n37255 & ~n37258 ;
  assign n37260 = n37259 ^ x508 ;
  assign n37261 = n37260 ^ x507 ;
  assign n37323 = n37262 ^ n37261 ;
  assign n37322 = n37320 & ~n37321 ;
  assign n37351 = n37323 ^ n37322 ;
  assign n37377 = n37351 ^ n36855 ;
  assign n37378 = n37377 ^ n37351 ;
  assign n37379 = n37378 ^ n37374 ;
  assign n37380 = n37376 & n37379 ;
  assign n37381 = n37380 ^ n37377 ;
  assign n37514 = n37381 ^ n36816 ;
  assign n37515 = n36245 & n37514 ;
  assign n37516 = n37515 ^ n36816 ;
  assign n37557 = n37516 ^ n35581 ;
  assign n37558 = n37557 ^ n37516 ;
  assign n37559 = n37558 ^ n37551 ;
  assign n37560 = ~n37556 & n37559 ;
  assign n37561 = n37560 ^ n37557 ;
  assign n37673 = n37561 ^ n35576 ;
  assign n37800 = n37673 ^ x193 ;
  assign n37702 = n37701 ^ n37675 ;
  assign n37703 = n37676 & ~n37702 ;
  assign n37704 = n37703 ^ x194 ;
  assign n37801 = n37800 ^ n37704 ;
  assign n37802 = n37799 & ~n37801 ;
  assign n37705 = n37704 ^ n37673 ;
  assign n37706 = n37704 ^ x193 ;
  assign n37707 = n37705 & n37706 ;
  assign n37708 = n37707 ^ x193 ;
  assign n37803 = n37708 ^ x192 ;
  assign n37517 = n37516 ^ n35576 ;
  assign n37562 = ~n37517 & ~n37561 ;
  assign n37563 = n37562 ^ n35576 ;
  assign n37263 = n37262 ^ n37260 ;
  assign n37264 = n37261 & n37263 ;
  assign n37265 = n37264 ^ x507 ;
  assign n37059 = n37058 ^ n35171 ;
  assign n37165 = n37059 & ~n37164 ;
  assign n37166 = n37165 ^ n35171 ;
  assign n37044 = n37043 ^ n37042 ;
  assign n37045 = n36573 ^ n36572 ;
  assign n37046 = n37045 ^ n36609 ;
  assign n37047 = n37046 ^ n37042 ;
  assign n37048 = n37047 ^ n37045 ;
  assign n37049 = ~n37044 & n37048 ;
  assign n37050 = n37049 ^ n37046 ;
  assign n37051 = n37050 ^ n36634 ;
  assign n37052 = ~n35984 & n37051 ;
  assign n37053 = n37052 ^ n36634 ;
  assign n37054 = n37053 ^ n35182 ;
  assign n37167 = n37166 ^ n37054 ;
  assign n37168 = n37167 ^ x506 ;
  assign n37325 = n37265 ^ n37168 ;
  assign n37324 = n37322 & n37323 ;
  assign n37384 = n37325 ^ n37324 ;
  assign n37509 = n37384 ^ n36812 ;
  assign n37352 = n37351 ^ n36816 ;
  assign n37382 = n37352 & ~n37381 ;
  assign n37383 = n37382 ^ n36816 ;
  assign n37510 = n37509 ^ n37383 ;
  assign n37511 = ~n36198 & ~n37510 ;
  assign n37512 = n37511 ^ n36812 ;
  assign n37513 = n37512 ^ n35571 ;
  assign n37671 = n37563 ^ n37513 ;
  assign n37804 = n37803 ^ n37671 ;
  assign n37805 = n37802 & n37804 ;
  assign n37385 = n37384 ^ n37383 ;
  assign n37269 = n37166 ^ n37053 ;
  assign n37272 = n37045 ^ n36634 ;
  assign n37273 = ~n37050 & ~n37272 ;
  assign n37274 = n37273 ^ n36634 ;
  assign n37270 = n36576 ^ n36574 ;
  assign n37271 = n37270 ^ n36650 ;
  assign n37275 = n37274 ^ n37271 ;
  assign n37276 = n36102 & n37275 ;
  assign n37277 = n37276 ^ n36650 ;
  assign n37278 = n37277 ^ n35182 ;
  assign n37279 = n37278 ^ n37166 ;
  assign n37280 = n37279 ^ n37277 ;
  assign n37281 = n37269 & n37280 ;
  assign n37282 = n37281 ^ n37278 ;
  assign n37283 = n37282 ^ n35375 ;
  assign n37347 = n37283 ^ x505 ;
  assign n37266 = n37265 ^ n37167 ;
  assign n37267 = n37168 & ~n37266 ;
  assign n37268 = n37267 ^ x506 ;
  assign n37348 = n37347 ^ n37268 ;
  assign n37326 = n37324 & ~n37325 ;
  assign n37349 = n37348 ^ n37326 ;
  assign n37386 = n37349 ^ n36812 ;
  assign n37387 = n37386 ^ n37349 ;
  assign n37388 = n37387 ^ n37383 ;
  assign n37389 = n37385 & n37388 ;
  assign n37390 = n37389 ^ n37386 ;
  assign n37567 = n37390 ^ n36867 ;
  assign n37568 = n36195 & ~n37567 ;
  assign n37569 = n37568 ^ n36867 ;
  assign n37712 = n37569 ^ n35566 ;
  assign n37564 = n37563 ^ n37512 ;
  assign n37565 = ~n37513 & n37564 ;
  assign n37566 = n37565 ^ n35571 ;
  assign n37713 = n37712 ^ n37566 ;
  assign n37806 = n37713 ^ x207 ;
  assign n37672 = n37671 ^ x192 ;
  assign n37709 = n37708 ^ n37671 ;
  assign n37710 = n37672 & ~n37709 ;
  assign n37711 = n37710 ^ x192 ;
  assign n37807 = n37806 ^ n37711 ;
  assign n37808 = ~n37805 & n37807 ;
  assign n37714 = n37713 ^ n37711 ;
  assign n37570 = n37569 ^ n37566 ;
  assign n37342 = n37277 ^ n35375 ;
  assign n37343 = n37282 & n37342 ;
  assign n37339 = n35467 ^ n35375 ;
  assign n37340 = n37339 ^ n36689 ;
  assign n37341 = n37340 ^ x504 ;
  assign n37344 = n37343 ^ n37341 ;
  assign n37335 = n37274 ^ n36650 ;
  assign n37336 = n37271 & n37335 ;
  assign n37332 = n36578 ^ n36577 ;
  assign n37333 = n37332 ^ n36689 ;
  assign n37334 = n37333 ^ n36650 ;
  assign n37337 = n37336 ^ n37334 ;
  assign n37338 = ~n36127 & n37337 ;
  assign n37345 = n37344 ^ n37338 ;
  assign n37284 = n37283 ^ n37268 ;
  assign n37327 = n37326 ^ n37268 ;
  assign n37330 = n37284 & n37327 ;
  assign n37285 = n37284 ^ n37268 ;
  assign n37328 = n37327 ^ n37285 ;
  assign n37329 = x505 & ~n37328 ;
  assign n37331 = n37330 ^ n37329 ;
  assign n37346 = n37345 ^ n37331 ;
  assign n37504 = n37346 ^ n36734 ;
  assign n37350 = n37349 ^ n36867 ;
  assign n37391 = ~n37350 & ~n37390 ;
  assign n37392 = n37391 ^ n36867 ;
  assign n37505 = n37504 ^ n37392 ;
  assign n37506 = ~n36190 & n37505 ;
  assign n37507 = n37506 ^ n36734 ;
  assign n37571 = n37507 ^ n35566 ;
  assign n37572 = n37571 ^ n37507 ;
  assign n37573 = n37572 ^ n37566 ;
  assign n37574 = ~n37570 & n37573 ;
  assign n37575 = n37574 ^ n37571 ;
  assign n37669 = n37575 ^ n35629 ;
  assign n37715 = n37669 ^ x207 ;
  assign n37716 = n37715 ^ n37669 ;
  assign n37717 = n37716 ^ n37711 ;
  assign n37718 = n37714 & n37717 ;
  assign n37719 = n37718 ^ n37715 ;
  assign n37809 = n37719 ^ x206 ;
  assign n37810 = n37808 & n37809 ;
  assign n37670 = n37669 ^ x206 ;
  assign n37720 = ~n37670 & n37719 ;
  assign n37721 = n37720 ^ x206 ;
  assign n37508 = n37507 ^ n35629 ;
  assign n37576 = n37508 & n37575 ;
  assign n37577 = n37576 ^ n35629 ;
  assign n37666 = n37577 ^ n35636 ;
  assign n37393 = n37392 ^ n37346 ;
  assign n37394 = n37392 ^ n36734 ;
  assign n37395 = ~n37393 & ~n37394 ;
  assign n37396 = n37395 ^ n36734 ;
  assign n37011 = n36909 ^ x487 ;
  assign n37012 = n37011 ^ n36805 ;
  assign n37500 = n37396 ^ n37012 ;
  assign n37501 = n36186 & ~n37500 ;
  assign n37502 = n37501 ^ n36805 ;
  assign n37667 = n37666 ^ n37502 ;
  assign n37668 = n37667 ^ x205 ;
  assign n37811 = n37721 ^ n37668 ;
  assign n37812 = ~n37810 & ~n37811 ;
  assign n37722 = n37721 ^ n37667 ;
  assign n37723 = ~n37668 & n37722 ;
  assign n37724 = n37723 ^ x205 ;
  assign n37813 = n37724 ^ x204 ;
  assign n37503 = n37502 ^ n35636 ;
  assign n37578 = n37577 ^ n37502 ;
  assign n37579 = ~n37503 & n37578 ;
  assign n37580 = n37579 ^ n35636 ;
  assign n37400 = n36910 ^ x486 ;
  assign n37401 = n37400 ^ n36907 ;
  assign n37495 = n37401 ^ n36886 ;
  assign n37397 = n37396 ^ n37011 ;
  assign n37398 = ~n37012 & ~n37397 ;
  assign n37399 = n37398 ^ n36805 ;
  assign n37496 = n37495 ^ n37399 ;
  assign n37497 = ~n36182 & ~n37496 ;
  assign n37498 = n37497 ^ n36886 ;
  assign n37499 = n37498 ^ n35563 ;
  assign n37664 = n37580 ^ n37499 ;
  assign n37814 = n37813 ^ n37664 ;
  assign n37815 = n37812 & n37814 ;
  assign n37665 = n37664 ^ x204 ;
  assign n37725 = n37724 ^ n37664 ;
  assign n37726 = n37665 & ~n37725 ;
  assign n37727 = n37726 ^ x204 ;
  assign n37816 = n37727 ^ x203 ;
  assign n37581 = n37580 ^ n37498 ;
  assign n37582 = n37499 & n37581 ;
  assign n37583 = n37582 ^ n35563 ;
  assign n37661 = n37583 ^ n35559 ;
  assign n37408 = n36916 ^ x485 ;
  assign n37402 = n37401 ^ n37399 ;
  assign n37403 = n36955 ^ n36886 ;
  assign n37404 = n37403 ^ n36955 ;
  assign n37405 = n37404 ^ n37399 ;
  assign n37406 = ~n37402 & n37405 ;
  assign n37407 = n37406 ^ n37403 ;
  assign n37491 = n37408 ^ n37407 ;
  assign n37492 = ~n36271 & n37491 ;
  assign n37493 = n37492 ^ n36955 ;
  assign n37662 = n37661 ^ n37493 ;
  assign n37817 = n37816 ^ n37662 ;
  assign n37818 = n37815 & n37817 ;
  assign n37663 = n37662 ^ x203 ;
  assign n37728 = n37727 ^ n37662 ;
  assign n37729 = n37663 & ~n37728 ;
  assign n37730 = n37729 ^ x203 ;
  assign n37819 = n37730 ^ x202 ;
  assign n37494 = n37493 ^ n35559 ;
  assign n37584 = n37583 ^ n37493 ;
  assign n37585 = ~n37494 & n37584 ;
  assign n37586 = n37585 ^ n35559 ;
  assign n37007 = n36903 ^ x484 ;
  assign n37008 = n37007 ^ n36918 ;
  assign n37410 = n37008 ^ n36955 ;
  assign n37409 = n37408 ^ n37008 ;
  assign n37411 = n37410 ^ n37409 ;
  assign n37412 = ~n37407 & ~n37411 ;
  assign n37413 = n37412 ^ n37410 ;
  assign n37487 = n37413 ^ n37009 ;
  assign n37488 = ~n36179 & n37487 ;
  assign n37489 = n37488 ^ n37009 ;
  assign n37490 = n37489 ^ n35555 ;
  assign n37659 = n37586 ^ n37490 ;
  assign n37820 = n37819 ^ n37659 ;
  assign n37821 = n37818 & n37820 ;
  assign n37660 = n37659 ^ x202 ;
  assign n37731 = n37730 ^ n37659 ;
  assign n37732 = n37660 & ~n37731 ;
  assign n37733 = n37732 ^ x202 ;
  assign n37822 = n37733 ^ x201 ;
  assign n37587 = n37586 ^ n37489 ;
  assign n37588 = ~n37490 & n37587 ;
  assign n37589 = n37588 ^ n35555 ;
  assign n37010 = n37009 ^ n37008 ;
  assign n37414 = n37010 & ~n37413 ;
  assign n37415 = n37414 ^ n37009 ;
  assign n37004 = n36922 ^ x483 ;
  assign n37005 = n37004 ^ n36901 ;
  assign n37006 = n37005 ^ n37003 ;
  assign n37483 = n37415 ^ n37006 ;
  assign n37484 = n36175 & n37483 ;
  assign n37485 = n37484 ^ n37003 ;
  assign n37486 = n37485 ^ n35653 ;
  assign n37734 = n37589 ^ n37486 ;
  assign n37823 = n37822 ^ n37734 ;
  assign n37824 = ~n37821 & ~n37823 ;
  assign n37735 = n37734 ^ n37733 ;
  assign n37590 = n37589 ^ n37485 ;
  assign n37591 = ~n37486 & ~n37590 ;
  assign n37592 = n37591 ^ n35653 ;
  assign n37416 = n37415 ^ n37003 ;
  assign n37417 = n37006 & n37416 ;
  assign n37418 = n37417 ^ n37005 ;
  assign n37002 = n37001 ^ n36965 ;
  assign n37479 = n37418 ^ n37002 ;
  assign n37480 = n36171 & ~n37479 ;
  assign n37481 = n37480 ^ n37001 ;
  assign n37482 = n37481 ^ n35551 ;
  assign n37736 = n37592 ^ n37482 ;
  assign n37737 = n37736 ^ x201 ;
  assign n37738 = n37737 ^ n37733 ;
  assign n37739 = n37738 ^ n37736 ;
  assign n37740 = ~n37735 & n37739 ;
  assign n37741 = n37740 ^ n37737 ;
  assign n37825 = n37741 ^ x200 ;
  assign n37826 = ~n37824 & ~n37825 ;
  assign n37419 = n37418 ^ n37001 ;
  assign n37420 = n37002 & ~n37419 ;
  assign n37421 = n37420 ^ n36965 ;
  assign n36999 = n36967 ^ n36965 ;
  assign n37000 = n36999 ^ n36998 ;
  assign n37597 = n37421 ^ n37000 ;
  assign n37598 = n36288 & n37597 ;
  assign n37599 = n37598 ^ n36998 ;
  assign n37593 = n37592 ^ n37481 ;
  assign n37594 = ~n37482 & n37593 ;
  assign n37595 = n37594 ^ n35551 ;
  assign n37596 = n37595 ^ n35547 ;
  assign n37657 = n37599 ^ n37596 ;
  assign n37743 = n37657 ^ x200 ;
  assign n37742 = n37736 ^ n37657 ;
  assign n37744 = n37743 ^ n37742 ;
  assign n37745 = n37741 & ~n37744 ;
  assign n37746 = n37745 ^ n37743 ;
  assign n37827 = n37746 ^ x215 ;
  assign n37828 = ~n37826 & ~n37827 ;
  assign n37422 = n37421 ^ n36998 ;
  assign n37423 = ~n37000 & ~n37422 ;
  assign n37424 = n37423 ^ n36999 ;
  assign n36995 = n36969 ^ n36968 ;
  assign n36997 = n36996 ^ n36995 ;
  assign n37476 = n37424 ^ n36997 ;
  assign n37477 = n36167 & n37476 ;
  assign n37478 = n37477 ^ n36996 ;
  assign n37655 = n37478 ^ n35542 ;
  assign n37600 = n37599 ^ n37595 ;
  assign n37601 = ~n37596 & n37600 ;
  assign n37602 = n37601 ^ n35547 ;
  assign n37656 = n37655 ^ n37602 ;
  assign n37789 = n37656 ^ x214 ;
  assign n37658 = n37657 ^ x215 ;
  assign n37747 = n37658 & ~n37746 ;
  assign n37748 = n37747 ^ x215 ;
  assign n37790 = n37789 ^ n37748 ;
  assign n37859 = n37828 ^ n37790 ;
  assign n37939 = n37859 ^ n37526 ;
  assign n37940 = n36581 & ~n37939 ;
  assign n37941 = n37940 ^ n37526 ;
  assign n37942 = ~n36209 & n37941 ;
  assign n37943 = n37942 ^ n36214 ;
  assign n37860 = ~n37526 & ~n37859 ;
  assign n37945 = n37860 ^ n37531 ;
  assign n37829 = n37790 & ~n37828 ;
  assign n37749 = n37748 ^ n37656 ;
  assign n37750 = n37748 ^ x214 ;
  assign n37751 = ~n37749 & n37750 ;
  assign n37752 = n37751 ^ x214 ;
  assign n37787 = n37752 ^ x213 ;
  assign n37603 = n37602 ^ n37478 ;
  assign n37604 = n37602 ^ n35542 ;
  assign n37605 = ~n37603 & ~n37604 ;
  assign n37606 = n37605 ^ n35542 ;
  assign n37753 = n37606 ^ n35538 ;
  assign n37427 = n36996 ^ n36992 ;
  assign n37425 = n37424 ^ n36995 ;
  assign n37426 = n36997 & n37425 ;
  assign n37428 = n37427 ^ n37426 ;
  assign n36993 = n36972 ^ n36970 ;
  assign n37472 = n37428 ^ n36993 ;
  assign n37473 = n36162 & n37472 ;
  assign n37474 = n37473 ^ n36992 ;
  assign n37754 = n37753 ^ n37474 ;
  assign n37788 = n37787 ^ n37754 ;
  assign n37858 = n37829 ^ n37788 ;
  assign n37946 = n37945 ^ n37858 ;
  assign n37947 = ~n36832 & ~n37946 ;
  assign n37944 = n37942 ^ n37531 ;
  assign n37948 = n37947 ^ n37944 ;
  assign n37949 = ~n37943 & n37948 ;
  assign n37950 = n37949 ^ n36214 ;
  assign n37861 = n37860 ^ n37858 ;
  assign n37830 = n37788 & n37829 ;
  assign n37755 = n37754 ^ n37752 ;
  assign n36994 = n36993 ^ n36992 ;
  assign n37429 = ~n36994 & n37428 ;
  assign n37430 = n37429 ^ n36993 ;
  assign n36990 = n36974 ^ n36973 ;
  assign n36991 = n36990 ^ n36989 ;
  assign n37469 = n37430 ^ n36991 ;
  assign n37470 = ~n36303 & ~n37469 ;
  assign n37471 = n37470 ^ n36989 ;
  assign n37652 = n37471 ^ n35534 ;
  assign n37475 = n37474 ^ n35538 ;
  assign n37607 = n37606 ^ n37474 ;
  assign n37608 = n37475 & ~n37607 ;
  assign n37609 = n37608 ^ n35538 ;
  assign n37653 = n37652 ^ n37609 ;
  assign n37756 = n37653 ^ x213 ;
  assign n37757 = n37756 ^ n37653 ;
  assign n37758 = n37757 ^ n37752 ;
  assign n37759 = ~n37755 & n37758 ;
  assign n37760 = n37759 ^ n37756 ;
  assign n37786 = n37760 ^ x212 ;
  assign n37856 = n37830 ^ n37786 ;
  assign n37862 = n37856 ^ n37531 ;
  assign n37863 = n37862 ^ n37858 ;
  assign n37864 = n37863 ^ n37856 ;
  assign n37865 = ~n37861 & n37864 ;
  assign n37866 = n37865 ^ n37862 ;
  assign n37935 = n37866 ^ n37523 ;
  assign n37936 = ~n36825 & n37935 ;
  assign n37937 = n37936 ^ n37523 ;
  assign n37938 = n37937 ^ n36205 ;
  assign n38033 = n37950 ^ n37938 ;
  assign n38025 = n37358 ^ n36580 ;
  assign n38026 = n38025 ^ n37940 ;
  assign n38027 = x423 & ~n38026 ;
  assign n38028 = n38027 ^ x422 ;
  assign n38029 = n37948 ^ n36214 ;
  assign n38030 = n38029 ^ n38027 ;
  assign n38031 = n38028 & ~n38030 ;
  assign n38032 = n38031 ^ x422 ;
  assign n38034 = n38033 ^ n38032 ;
  assign n38104 = n38034 ^ x421 ;
  assign n38105 = n38026 ^ x423 ;
  assign n38106 = n38029 ^ n38028 ;
  assign n38107 = ~n38105 & n38106 ;
  assign n38108 = n38104 & n38107 ;
  assign n38035 = n38032 ^ x421 ;
  assign n38036 = ~n38034 & n38035 ;
  assign n38037 = n38036 ^ x421 ;
  assign n37951 = n37950 ^ n37937 ;
  assign n37952 = ~n37938 & ~n37951 ;
  assign n37953 = n37952 ^ n36205 ;
  assign n37857 = n37856 ^ n37523 ;
  assign n37867 = ~n37857 & n37866 ;
  assign n37868 = n37867 ^ n37523 ;
  assign n37930 = n37868 ^ n37518 ;
  assign n37433 = n36990 ^ n36986 ;
  assign n37431 = n37430 ^ n36989 ;
  assign n37432 = n36991 & n37431 ;
  assign n37434 = n37433 ^ n37432 ;
  assign n36987 = n36976 ^ n36975 ;
  assign n37614 = n37434 ^ n36987 ;
  assign n37615 = n36158 & ~n37614 ;
  assign n37616 = n37615 ^ n36986 ;
  assign n37763 = n37616 ^ n35677 ;
  assign n37610 = n37609 ^ n37471 ;
  assign n37611 = n37609 ^ n35534 ;
  assign n37612 = ~n37610 & ~n37611 ;
  assign n37613 = n37612 ^ n35534 ;
  assign n37764 = n37763 ^ n37613 ;
  assign n37832 = n37764 ^ x211 ;
  assign n37654 = n37653 ^ x212 ;
  assign n37761 = ~n37654 & n37760 ;
  assign n37762 = n37761 ^ x212 ;
  assign n37833 = n37832 ^ n37762 ;
  assign n37831 = ~n37786 & n37830 ;
  assign n37854 = n37833 ^ n37831 ;
  assign n37931 = n37930 ^ n37854 ;
  assign n37932 = ~n36839 & n37931 ;
  assign n37933 = n37932 ^ n37518 ;
  assign n37934 = n37933 ^ n36203 ;
  assign n38023 = n37953 ^ n37934 ;
  assign n38024 = n38023 ^ x420 ;
  assign n38109 = n38037 ^ n38024 ;
  assign n38110 = n38108 & ~n38109 ;
  assign n37954 = n37953 ^ n37933 ;
  assign n37955 = ~n37934 & n37954 ;
  assign n37956 = n37955 ^ n36203 ;
  assign n38042 = n37956 ^ n36230 ;
  assign n37855 = n37854 ^ n37518 ;
  assign n37869 = n37868 ^ n37854 ;
  assign n37870 = ~n37855 & n37869 ;
  assign n37871 = n37870 ^ n37518 ;
  assign n37765 = n37764 ^ n37762 ;
  assign n37617 = n37616 ^ n37613 ;
  assign n37620 = n37613 ^ n35677 ;
  assign n37621 = n37617 & ~n37620 ;
  assign n36988 = n36987 ^ n36986 ;
  assign n37435 = ~n36988 & ~n37434 ;
  assign n37436 = n37435 ^ n36987 ;
  assign n36984 = n36979 ^ n36977 ;
  assign n36985 = n36984 ^ n36983 ;
  assign n37465 = n37436 ^ n36985 ;
  assign n37466 = n36154 & ~n37465 ;
  assign n37467 = n37466 ^ n36983 ;
  assign n37618 = n37467 ^ n35677 ;
  assign n37622 = n37621 ^ n37618 ;
  assign n37650 = n37622 ^ n35508 ;
  assign n37766 = n37650 ^ x211 ;
  assign n37767 = n37766 ^ n37762 ;
  assign n37768 = n37767 ^ n37650 ;
  assign n37769 = n37765 & n37768 ;
  assign n37770 = n37769 ^ n37766 ;
  assign n37835 = n37770 ^ x210 ;
  assign n37834 = n37831 & ~n37833 ;
  assign n37852 = n37835 ^ n37834 ;
  assign n37853 = n37852 ^ n37546 ;
  assign n37957 = n37871 ^ n37853 ;
  assign n37958 = ~n36820 & n37957 ;
  assign n37959 = n37958 ^ n37546 ;
  assign n38043 = n38042 ^ n37959 ;
  assign n38038 = n38037 ^ n38023 ;
  assign n38039 = ~n38024 & n38038 ;
  assign n38040 = n38039 ^ x420 ;
  assign n38041 = n38040 ^ x419 ;
  assign n38111 = n38043 ^ n38041 ;
  assign n38112 = n38110 & n38111 ;
  assign n37960 = n37959 ^ n37956 ;
  assign n37961 = n37959 ^ n36230 ;
  assign n37962 = n37960 & n37961 ;
  assign n37963 = n37962 ^ n36230 ;
  assign n38021 = n37963 ^ n36237 ;
  assign n37872 = n37871 ^ n37852 ;
  assign n37873 = ~n37853 & n37872 ;
  assign n37874 = n37873 ^ n37546 ;
  assign n37439 = n36984 ^ n36804 ;
  assign n37437 = n37436 ^ n36983 ;
  assign n37438 = n36985 & n37437 ;
  assign n37440 = n37439 ^ n37438 ;
  assign n36981 = n36980 ^ n36964 ;
  assign n37625 = n37440 ^ n36981 ;
  assign n37626 = ~n36150 & ~n37625 ;
  assign n37627 = n37626 ^ n36804 ;
  assign n37648 = n37627 ^ n35529 ;
  assign n37468 = n37467 ^ n35508 ;
  assign n37623 = ~n37468 & ~n37622 ;
  assign n37624 = n37623 ^ n35508 ;
  assign n37649 = n37648 ^ n37624 ;
  assign n37837 = n37649 ^ x209 ;
  assign n37651 = n37650 ^ x210 ;
  assign n37771 = ~n37651 & n37770 ;
  assign n37772 = n37771 ^ x210 ;
  assign n37838 = n37837 ^ n37772 ;
  assign n37836 = n37834 & ~n37835 ;
  assign n37850 = n37838 ^ n37836 ;
  assign n37851 = n37850 ^ n37553 ;
  assign n37926 = n37874 ^ n37851 ;
  assign n37927 = ~n36855 & n37926 ;
  assign n37928 = n37927 ^ n37553 ;
  assign n38022 = n38021 ^ n37928 ;
  assign n38113 = n38022 ^ x418 ;
  assign n38044 = n38043 ^ n38040 ;
  assign n38045 = n38041 & ~n38044 ;
  assign n38046 = n38045 ^ x419 ;
  assign n38114 = n38113 ^ n38046 ;
  assign n38115 = ~n38112 & ~n38114 ;
  assign n38047 = n38046 ^ n38022 ;
  assign n38048 = n38046 ^ x418 ;
  assign n38049 = ~n38047 & n38048 ;
  assign n38050 = n38049 ^ x418 ;
  assign n37929 = n37928 ^ n36237 ;
  assign n37964 = n37963 ^ n37928 ;
  assign n37965 = ~n37929 & ~n37964 ;
  assign n37966 = n37965 ^ n36237 ;
  assign n37875 = n37874 ^ n37850 ;
  assign n37876 = ~n37851 & n37875 ;
  assign n37877 = n37876 ^ n37553 ;
  assign n37773 = n37772 ^ n37649 ;
  assign n37774 = n37772 ^ x209 ;
  assign n37775 = n37773 & n37774 ;
  assign n37776 = n37775 ^ x209 ;
  assign n37628 = n37627 ^ n37624 ;
  assign n37444 = n37289 ^ n37288 ;
  assign n37460 = n37444 ^ n37072 ;
  assign n36982 = n36981 ^ n36804 ;
  assign n37441 = ~n36982 & n37440 ;
  assign n37442 = n37441 ^ n36981 ;
  assign n37461 = n37460 ^ n37442 ;
  assign n37462 = n36325 & n37461 ;
  assign n37463 = n37462 ^ n37072 ;
  assign n37629 = n37463 ^ n35529 ;
  assign n37630 = n37629 ^ n37624 ;
  assign n37631 = n37630 ^ n37463 ;
  assign n37632 = ~n37628 & n37631 ;
  assign n37633 = n37632 ^ n37629 ;
  assign n37646 = n37633 ^ n35526 ;
  assign n37647 = n37646 ^ x208 ;
  assign n37840 = n37776 ^ n37647 ;
  assign n37839 = n37836 & ~n37838 ;
  assign n37848 = n37840 ^ n37839 ;
  assign n37849 = n37848 ^ n37514 ;
  assign n37922 = n37877 ^ n37849 ;
  assign n37923 = ~n36816 & n37922 ;
  assign n37924 = n37923 ^ n37514 ;
  assign n37925 = n37924 ^ n36245 ;
  assign n38019 = n37966 ^ n37925 ;
  assign n38020 = n38019 ^ x417 ;
  assign n38116 = n38050 ^ n38020 ;
  assign n38117 = ~n38115 & n38116 ;
  assign n38051 = n38050 ^ n38019 ;
  assign n38052 = n38020 & ~n38051 ;
  assign n38053 = n38052 ^ x417 ;
  assign n38118 = n38053 ^ x416 ;
  assign n37967 = n37966 ^ n37924 ;
  assign n37968 = n37925 & ~n37967 ;
  assign n37969 = n37968 ^ n36245 ;
  assign n37878 = n37877 ^ n37848 ;
  assign n37879 = ~n37849 & ~n37878 ;
  assign n37880 = n37879 ^ n37514 ;
  assign n37917 = n37880 ^ n37510 ;
  assign n37451 = n37292 ^ n37290 ;
  assign n37443 = n37442 ^ n37072 ;
  assign n37447 = n37444 ^ n37442 ;
  assign n37448 = ~n37443 & n37447 ;
  assign n37445 = n37444 ^ n37068 ;
  assign n37449 = n37448 ^ n37445 ;
  assign n37637 = n37451 ^ n37449 ;
  assign n37638 = n36334 & n37637 ;
  assign n37639 = n37638 ^ n37068 ;
  assign n37464 = n37463 ^ n35526 ;
  assign n37634 = ~n37464 & n37633 ;
  assign n37635 = n37634 ^ n35526 ;
  assign n37636 = n37635 ^ n35827 ;
  assign n37781 = n37639 ^ n37636 ;
  assign n37777 = n37776 ^ n37646 ;
  assign n37778 = n37647 & ~n37777 ;
  assign n37779 = n37778 ^ x208 ;
  assign n37780 = n37779 ^ x223 ;
  assign n37842 = n37781 ^ n37780 ;
  assign n37841 = n37839 & n37840 ;
  assign n37846 = n37842 ^ n37841 ;
  assign n37918 = n37917 ^ n37846 ;
  assign n37919 = ~n36812 & ~n37918 ;
  assign n37920 = n37919 ^ n37510 ;
  assign n37921 = n37920 ^ n36198 ;
  assign n38017 = n37969 ^ n37921 ;
  assign n38119 = n38118 ^ n38017 ;
  assign n38120 = ~n38117 & ~n38119 ;
  assign n38018 = n38017 ^ x416 ;
  assign n38054 = n38053 ^ n38017 ;
  assign n38055 = n38018 & ~n38054 ;
  assign n38056 = n38055 ^ x416 ;
  assign n38121 = n38056 ^ x431 ;
  assign n37970 = n37969 ^ n37920 ;
  assign n37971 = n37921 & n37970 ;
  assign n37972 = n37971 ^ n36198 ;
  assign n37847 = n37846 ^ n37510 ;
  assign n37881 = n37880 ^ n37846 ;
  assign n37882 = ~n37847 & ~n37881 ;
  assign n37883 = n37882 ^ n37510 ;
  assign n37843 = ~n37841 & ~n37842 ;
  assign n37782 = n37781 ^ n37779 ;
  assign n37783 = n37780 & ~n37782 ;
  assign n37784 = n37783 ^ x223 ;
  assign n37640 = n37639 ^ n37635 ;
  assign n37641 = n37636 & n37640 ;
  assign n37642 = n37641 ^ n35827 ;
  assign n37643 = n37642 ^ n35905 ;
  assign n37450 = n37295 ^ n37293 ;
  assign n37453 = n37450 ^ n37068 ;
  assign n37452 = n37451 ^ n37450 ;
  assign n37454 = n37453 ^ n37452 ;
  assign n37455 = n37449 & n37454 ;
  assign n37456 = n37455 ^ n37453 ;
  assign n37457 = n37456 ^ n37064 ;
  assign n37458 = ~n36347 & ~n37457 ;
  assign n37459 = n37458 ^ n37064 ;
  assign n37644 = n37643 ^ n37459 ;
  assign n37645 = n37644 ^ x222 ;
  assign n37785 = n37784 ^ n37645 ;
  assign n37844 = n37843 ^ n37785 ;
  assign n37845 = n37844 ^ n37567 ;
  assign n37913 = n37883 ^ n37845 ;
  assign n37914 = n36867 & n37913 ;
  assign n37915 = n37914 ^ n37567 ;
  assign n37916 = n37915 ^ n36195 ;
  assign n38015 = n37972 ^ n37916 ;
  assign n38122 = n38121 ^ n38015 ;
  assign n38123 = n38120 & ~n38122 ;
  assign n38016 = n38015 ^ x431 ;
  assign n38057 = n38056 ^ n38015 ;
  assign n38058 = n38016 & ~n38057 ;
  assign n38059 = n38058 ^ x431 ;
  assign n38124 = n38059 ^ x430 ;
  assign n37973 = n37972 ^ n37915 ;
  assign n37974 = ~n37916 & ~n37973 ;
  assign n37975 = n37974 ^ n36195 ;
  assign n38012 = n37975 ^ n36190 ;
  assign n37906 = n37785 & n37843 ;
  assign n37900 = n37784 ^ n37644 ;
  assign n37901 = n37784 ^ x222 ;
  assign n37902 = n37900 & n37901 ;
  assign n37903 = n37902 ^ x222 ;
  assign n37904 = n37903 ^ x221 ;
  assign n37896 = n37642 ^ n37459 ;
  assign n37897 = ~n37643 & n37896 ;
  assign n37898 = n37897 ^ n35905 ;
  assign n37889 = n37450 ^ n37064 ;
  assign n37890 = n37456 & ~n37889 ;
  assign n37891 = n37890 ^ n37064 ;
  assign n37887 = n37298 ^ n37296 ;
  assign n37888 = n37887 ^ n37060 ;
  assign n37892 = n37891 ^ n37888 ;
  assign n37893 = ~n36509 & ~n37892 ;
  assign n37894 = n37893 ^ n37060 ;
  assign n37895 = n37894 ^ n35929 ;
  assign n37899 = n37898 ^ n37895 ;
  assign n37905 = n37904 ^ n37899 ;
  assign n37907 = n37906 ^ n37905 ;
  assign n37908 = n37907 ^ n37505 ;
  assign n37884 = n37883 ^ n37844 ;
  assign n37885 = ~n37845 & n37884 ;
  assign n37886 = n37885 ^ n37567 ;
  assign n37909 = n37908 ^ n37886 ;
  assign n37910 = ~n36734 & n37909 ;
  assign n37911 = n37910 ^ n37505 ;
  assign n38013 = n38012 ^ n37911 ;
  assign n38125 = n38124 ^ n38013 ;
  assign n38126 = ~n38123 & ~n38125 ;
  assign n38014 = n38013 ^ x430 ;
  assign n38060 = n38059 ^ n38013 ;
  assign n38061 = ~n38014 & n38060 ;
  assign n38062 = n38061 ^ x430 ;
  assign n38127 = n38062 ^ x429 ;
  assign n38004 = ~n37905 & ~n37906 ;
  assign n37999 = n37899 ^ x221 ;
  assign n38000 = n37903 ^ n37899 ;
  assign n38001 = ~n37999 & n38000 ;
  assign n38002 = n38001 ^ x221 ;
  assign n37992 = n37898 ^ n37894 ;
  assign n37993 = n37898 ^ n35929 ;
  assign n37994 = n37992 & n37993 ;
  assign n37995 = n37994 ^ n35929 ;
  assign n37996 = n37995 ^ n35948 ;
  assign n37988 = n37300 ^ n37299 ;
  assign n37986 = n37156 ^ n37060 ;
  assign n37983 = n37891 ^ n37887 ;
  assign n37984 = n37891 ^ n37060 ;
  assign n37985 = ~n37983 & ~n37984 ;
  assign n37987 = n37986 ^ n37985 ;
  assign n37989 = n37988 ^ n37987 ;
  assign n37990 = n36591 & n37989 ;
  assign n37991 = n37990 ^ n37156 ;
  assign n37997 = n37996 ^ n37991 ;
  assign n37998 = n37997 ^ x220 ;
  assign n38003 = n38002 ^ n37998 ;
  assign n38005 = n38004 ^ n38003 ;
  assign n37979 = n37907 ^ n37886 ;
  assign n37980 = ~n37908 & ~n37979 ;
  assign n37981 = n37980 ^ n37505 ;
  assign n37982 = n37981 ^ n37500 ;
  assign n38006 = n38005 ^ n37982 ;
  assign n38007 = n36805 & ~n38006 ;
  assign n38008 = n38007 ^ n37500 ;
  assign n38009 = n38008 ^ n36186 ;
  assign n37912 = n37911 ^ n36190 ;
  assign n37976 = n37975 ^ n37911 ;
  assign n37977 = ~n37912 & ~n37976 ;
  assign n37978 = n37977 ^ n36190 ;
  assign n38010 = n38009 ^ n37978 ;
  assign n38128 = n38127 ^ n38010 ;
  assign n38129 = n38126 & n38128 ;
  assign n38094 = ~n38003 & n38004 ;
  assign n38088 = n38002 ^ n37997 ;
  assign n38089 = n38002 ^ x220 ;
  assign n38090 = n38088 & n38089 ;
  assign n38091 = n38090 ^ x220 ;
  assign n38092 = n38091 ^ x219 ;
  assign n38073 = n37995 ^ n37991 ;
  assign n38076 = n37988 ^ n37156 ;
  assign n38077 = ~n37987 & ~n38076 ;
  assign n38078 = n38077 ^ n37156 ;
  assign n38074 = n37301 ^ n37286 ;
  assign n38075 = n38074 ^ n37056 ;
  assign n38079 = n38078 ^ n38075 ;
  assign n38080 = n36609 & ~n38079 ;
  assign n38081 = n38080 ^ n37056 ;
  assign n38082 = n38081 ^ n35948 ;
  assign n38083 = n38082 ^ n38081 ;
  assign n38084 = n38083 ^ n37995 ;
  assign n38085 = ~n38073 & ~n38084 ;
  assign n38086 = n38085 ^ n38082 ;
  assign n38087 = n38086 ^ n35965 ;
  assign n38093 = n38092 ^ n38087 ;
  assign n38095 = n38094 ^ n38093 ;
  assign n38096 = n38095 ^ n37496 ;
  assign n38069 = n38005 ^ n37500 ;
  assign n38070 = n38005 ^ n37981 ;
  assign n38071 = ~n38069 & ~n38070 ;
  assign n38072 = n38071 ^ n37500 ;
  assign n38097 = n38096 ^ n38072 ;
  assign n38098 = n36886 & ~n38097 ;
  assign n38099 = n38098 ^ n37496 ;
  assign n38100 = n38099 ^ n36182 ;
  assign n38066 = n38008 ^ n37978 ;
  assign n38067 = ~n38009 & ~n38066 ;
  assign n38068 = n38067 ^ n36186 ;
  assign n38101 = n38100 ^ n38068 ;
  assign n38102 = n38101 ^ x428 ;
  assign n38011 = n38010 ^ x429 ;
  assign n38063 = n38062 ^ n38010 ;
  assign n38064 = n38011 & ~n38063 ;
  assign n38065 = n38064 ^ x429 ;
  assign n38103 = n38102 ^ n38065 ;
  assign n38130 = n38129 ^ n38103 ;
  assign n38131 = n38130 ^ n37859 ;
  assign n39277 = n38131 ^ n37526 ;
  assign n38132 = n37859 ^ n36581 ;
  assign n38133 = n38132 ^ n37358 ;
  assign n38134 = n38133 ^ n38130 ;
  assign n38135 = n38131 & n38134 ;
  assign n38136 = n38135 ^ n38132 ;
  assign n38187 = x135 & n38136 ;
  assign n38188 = n38187 ^ x134 ;
  assign n38181 = n37939 & n38130 ;
  assign n38182 = n38181 ^ n37946 ;
  assign n38179 = n38103 & n38129 ;
  assign n38170 = n38093 & n38094 ;
  assign n38165 = n38087 ^ x219 ;
  assign n38166 = n38091 ^ n38087 ;
  assign n38167 = n38165 & ~n38166 ;
  assign n38168 = n38167 ^ x219 ;
  assign n38153 = n37303 ^ n37302 ;
  assign n38154 = n38153 ^ n37051 ;
  assign n38149 = n38078 ^ n38074 ;
  assign n38150 = n38078 ^ n37056 ;
  assign n38151 = ~n38149 & ~n38150 ;
  assign n38152 = n38151 ^ n37056 ;
  assign n38155 = n38154 ^ n38152 ;
  assign n38156 = ~n36634 & n38155 ;
  assign n38157 = n38156 ^ n37051 ;
  assign n38159 = n38157 ^ n35965 ;
  assign n38158 = n38157 ^ n38081 ;
  assign n38160 = n38159 ^ n38158 ;
  assign n38161 = ~n38086 & ~n38160 ;
  assign n38162 = n38161 ^ n38159 ;
  assign n38163 = n38162 ^ n35984 ;
  assign n38164 = n38163 ^ x218 ;
  assign n38169 = n38168 ^ n38164 ;
  assign n38171 = n38170 ^ n38169 ;
  assign n38172 = n38171 ^ n37491 ;
  assign n38146 = n38095 ^ n38072 ;
  assign n38147 = n38096 & ~n38146 ;
  assign n38148 = n38147 ^ n37496 ;
  assign n38173 = n38172 ^ n38148 ;
  assign n38174 = ~n36955 & n38173 ;
  assign n38175 = n38174 ^ n37491 ;
  assign n38142 = n38099 ^ n38068 ;
  assign n38143 = n38100 & n38142 ;
  assign n38144 = n38143 ^ n36182 ;
  assign n38145 = n38144 ^ n36271 ;
  assign n38176 = n38175 ^ n38145 ;
  assign n38177 = n38176 ^ x427 ;
  assign n38139 = n38101 ^ n38065 ;
  assign n38140 = n38102 & ~n38139 ;
  assign n38141 = n38140 ^ x428 ;
  assign n38178 = n38177 ^ n38141 ;
  assign n38180 = n38179 ^ n38178 ;
  assign n38183 = n38182 ^ n38180 ;
  assign n38184 = n37531 & n38183 ;
  assign n38137 = n36581 & ~n38136 ;
  assign n38138 = n38137 ^ n37946 ;
  assign n38185 = n38184 ^ n38138 ;
  assign n38186 = n38185 ^ n36832 ;
  assign n38189 = n38188 ^ n38186 ;
  assign n38223 = n38169 & ~n38170 ;
  assign n38210 = n38153 ^ n38152 ;
  assign n38211 = n37305 ^ n37304 ;
  assign n38212 = n38211 ^ n37051 ;
  assign n38213 = n38212 ^ n38211 ;
  assign n38214 = n38213 ^ n38152 ;
  assign n38215 = ~n38210 & ~n38214 ;
  assign n38216 = n38215 ^ n38212 ;
  assign n38217 = n38216 ^ n37275 ;
  assign n38218 = ~n36650 & n38217 ;
  assign n38219 = n38218 ^ n37275 ;
  assign n38206 = n38157 ^ n35984 ;
  assign n38207 = ~n38162 & ~n38206 ;
  assign n38208 = n38207 ^ n35984 ;
  assign n38209 = n38208 ^ n36102 ;
  assign n38220 = n38219 ^ n38209 ;
  assign n38221 = n38220 ^ x217 ;
  assign n38202 = n38168 ^ n38163 ;
  assign n38203 = n38168 ^ x218 ;
  assign n38204 = n38202 & n38203 ;
  assign n38205 = n38204 ^ x218 ;
  assign n38222 = n38221 ^ n38205 ;
  assign n38224 = n38223 ^ n38222 ;
  assign n38225 = n38224 ^ n37487 ;
  assign n38199 = n38171 ^ n38148 ;
  assign n38200 = ~n38172 & ~n38199 ;
  assign n38201 = n38200 ^ n37491 ;
  assign n38226 = n38225 ^ n38201 ;
  assign n38227 = ~n37009 & ~n38226 ;
  assign n38228 = n38227 ^ n37487 ;
  assign n38194 = n38175 ^ n36271 ;
  assign n38195 = n38175 ^ n38144 ;
  assign n38196 = ~n38194 & n38195 ;
  assign n38197 = n38196 ^ n36271 ;
  assign n38198 = n38197 ^ n36179 ;
  assign n38229 = n38228 ^ n38198 ;
  assign n38230 = n38229 ^ x426 ;
  assign n38191 = n38176 ^ n38141 ;
  assign n38192 = n38177 & ~n38191 ;
  assign n38193 = n38192 ^ x427 ;
  assign n38231 = n38230 ^ n38193 ;
  assign n38190 = ~n38178 & ~n38179 ;
  assign n38295 = n38231 ^ n38190 ;
  assign n38825 = n38295 ^ n37935 ;
  assign n38296 = n38181 ^ n38180 ;
  assign n38297 = n38182 & n38296 ;
  assign n38298 = n38297 ^ n37946 ;
  assign n38826 = n38825 ^ n38298 ;
  assign n38827 = n37523 & ~n38826 ;
  assign n38828 = n38827 ^ n37935 ;
  assign n39037 = n38828 ^ n36825 ;
  assign n38829 = n38137 ^ n36832 ;
  assign n38830 = n38185 & ~n38829 ;
  assign n38831 = n38830 ^ n36832 ;
  assign n39038 = n39037 ^ n38831 ;
  assign n39033 = n38187 ^ n38186 ;
  assign n39034 = n38188 & ~n39033 ;
  assign n39035 = n39034 ^ x134 ;
  assign n39039 = n39038 ^ n39035 ;
  assign n39215 = n39039 ^ x133 ;
  assign n39216 = n38189 & n39215 ;
  assign n39036 = n39035 ^ x133 ;
  assign n39040 = n39036 & ~n39039 ;
  assign n39041 = n39040 ^ x133 ;
  assign n38299 = n38298 ^ n38295 ;
  assign n38300 = n38298 ^ n37935 ;
  assign n38301 = n38299 & ~n38300 ;
  assign n38302 = n38301 ^ n37935 ;
  assign n38261 = n38224 ^ n38201 ;
  assign n38262 = ~n38225 & n38261 ;
  assign n38263 = n38262 ^ n37487 ;
  assign n38264 = n38263 ^ n37483 ;
  assign n38259 = ~n38222 & ~n38223 ;
  assign n38255 = n38220 ^ n38205 ;
  assign n38256 = ~n38221 & n38255 ;
  assign n38253 = x217 ^ x216 ;
  assign n38248 = n38211 ^ n37275 ;
  assign n38249 = n38216 & n38248 ;
  assign n38245 = n37308 ^ n37306 ;
  assign n38246 = n38245 ^ n37337 ;
  assign n38247 = n38246 ^ n38211 ;
  assign n38250 = n38249 ^ n38247 ;
  assign n38251 = ~n36689 & ~n38250 ;
  assign n38243 = n36127 ^ n36102 ;
  assign n38244 = n38243 ^ n37337 ;
  assign n38252 = n38251 ^ n38244 ;
  assign n38254 = n38253 ^ n38252 ;
  assign n38257 = n38256 ^ n38254 ;
  assign n38240 = n38219 ^ n38208 ;
  assign n38241 = n38219 ^ n36102 ;
  assign n38242 = n38240 & n38241 ;
  assign n38258 = n38257 ^ n38242 ;
  assign n38260 = n38259 ^ n38258 ;
  assign n38265 = n38264 ^ n38260 ;
  assign n38266 = n37003 & ~n38265 ;
  assign n38267 = n38266 ^ n37483 ;
  assign n38268 = n38267 ^ n36175 ;
  assign n38236 = n38228 ^ n36179 ;
  assign n38237 = n38228 ^ n38197 ;
  assign n38238 = ~n38236 & n38237 ;
  assign n38239 = n38238 ^ n36179 ;
  assign n38269 = n38268 ^ n38239 ;
  assign n38270 = n38269 ^ x425 ;
  assign n38233 = n38229 ^ n38193 ;
  assign n38234 = n38230 & ~n38233 ;
  assign n38235 = n38234 ^ x426 ;
  assign n38271 = n38270 ^ n38235 ;
  assign n38232 = ~n38190 & n38231 ;
  assign n38293 = n38271 ^ n38232 ;
  assign n38294 = n38293 ^ n37931 ;
  assign n38836 = n38302 ^ n38294 ;
  assign n38837 = n37518 & n38836 ;
  assign n38838 = n38837 ^ n37931 ;
  assign n39030 = n38838 ^ n36839 ;
  assign n38832 = n38831 ^ n38828 ;
  assign n38833 = n38831 ^ n36825 ;
  assign n38834 = n38832 & n38833 ;
  assign n38835 = n38834 ^ n36825 ;
  assign n39031 = n39030 ^ n38835 ;
  assign n39032 = n39031 ^ x132 ;
  assign n39217 = n39041 ^ n39032 ;
  assign n39218 = n39216 & n39217 ;
  assign n38839 = n38838 ^ n38835 ;
  assign n38303 = n38302 ^ n38293 ;
  assign n38304 = n38294 & ~n38303 ;
  assign n38305 = n38304 ^ n37931 ;
  assign n38820 = n38305 ^ n37957 ;
  assign n38287 = n38269 ^ n38235 ;
  assign n38288 = ~n38270 & n38287 ;
  assign n38289 = n38288 ^ x425 ;
  assign n38282 = n38267 ^ n38239 ;
  assign n38283 = n38268 & n38282 ;
  assign n38284 = n38283 ^ n36175 ;
  assign n38275 = n38263 ^ n38260 ;
  assign n38276 = n38264 & n38275 ;
  assign n38277 = n38276 ^ n37483 ;
  assign n38273 = n37685 ^ x199 ;
  assign n38274 = n38273 ^ n37479 ;
  assign n38278 = n38277 ^ n38274 ;
  assign n38279 = n37001 & ~n38278 ;
  assign n38280 = n38279 ^ n37479 ;
  assign n38281 = n38280 ^ n36171 ;
  assign n38285 = n38284 ^ n38281 ;
  assign n38286 = n38285 ^ x424 ;
  assign n38290 = n38289 ^ n38286 ;
  assign n38272 = n38232 & ~n38271 ;
  assign n38291 = n38290 ^ n38272 ;
  assign n38821 = n38820 ^ n38291 ;
  assign n38822 = n37546 & n38821 ;
  assign n38823 = n38822 ^ n37957 ;
  assign n38840 = n38823 ^ n36839 ;
  assign n38841 = n38840 ^ n38823 ;
  assign n38842 = n38841 ^ n38835 ;
  assign n38843 = n38839 & n38842 ;
  assign n38844 = n38843 ^ n38840 ;
  assign n39029 = n38844 ^ n36820 ;
  assign n39219 = n39029 ^ x131 ;
  assign n39042 = n39041 ^ n39031 ;
  assign n39043 = n39032 & ~n39042 ;
  assign n39044 = n39043 ^ x132 ;
  assign n39220 = n39219 ^ n39044 ;
  assign n39221 = n39218 & n39220 ;
  assign n38311 = n38289 ^ n38285 ;
  assign n38320 = n37686 ^ x198 ;
  assign n38321 = n38320 ^ n37683 ;
  assign n38322 = n38321 ^ n37597 ;
  assign n38316 = n38277 ^ n37479 ;
  assign n38317 = n38277 ^ n38273 ;
  assign n38318 = ~n38316 & ~n38317 ;
  assign n38319 = n38318 ^ n37479 ;
  assign n38323 = n38322 ^ n38319 ;
  assign n38324 = n36998 & ~n38323 ;
  assign n38325 = n38324 ^ n37597 ;
  assign n38312 = n38284 ^ n38280 ;
  assign n38313 = ~n38281 & n38312 ;
  assign n38314 = n38313 ^ n36171 ;
  assign n38315 = n38314 ^ n36288 ;
  assign n38326 = n38325 ^ n38315 ;
  assign n38327 = n38326 ^ x424 ;
  assign n38328 = n38327 ^ n38326 ;
  assign n38329 = n38328 ^ n38289 ;
  assign n38330 = n38311 & n38329 ;
  assign n38331 = n38330 ^ n38327 ;
  assign n38332 = n38331 ^ x439 ;
  assign n38310 = n38272 & ~n38290 ;
  assign n38333 = n38332 ^ n38310 ;
  assign n38292 = n38291 ^ n37957 ;
  assign n38306 = n38305 ^ n38291 ;
  assign n38307 = n38292 & ~n38306 ;
  assign n38308 = n38307 ^ n37957 ;
  assign n38334 = n38333 ^ n38308 ;
  assign n38817 = n38334 ^ n37926 ;
  assign n38818 = n37553 & ~n38817 ;
  assign n38819 = n38818 ^ n37926 ;
  assign n39049 = n38819 ^ n36855 ;
  assign n38824 = n38823 ^ n36820 ;
  assign n38845 = ~n38824 & n38844 ;
  assign n38846 = n38845 ^ n36820 ;
  assign n39050 = n39049 ^ n38846 ;
  assign n39052 = n39050 ^ x130 ;
  assign n39045 = n39044 ^ n39029 ;
  assign n39046 = n39044 ^ x131 ;
  assign n39047 = ~n39045 & n39046 ;
  assign n39048 = n39047 ^ x131 ;
  assign n39222 = n39052 ^ n39048 ;
  assign n39223 = n39221 & n39222 ;
  assign n38847 = n38846 ^ n38819 ;
  assign n38354 = n38326 ^ x439 ;
  assign n38355 = ~n38331 & n38354 ;
  assign n38356 = n38355 ^ x439 ;
  assign n38339 = n38325 ^ n38314 ;
  assign n38343 = n37791 ^ n37476 ;
  assign n38340 = n38321 ^ n38319 ;
  assign n38341 = n38322 & n38340 ;
  assign n38342 = n38341 ^ n37597 ;
  assign n38344 = n38343 ^ n38342 ;
  assign n38345 = n36996 & ~n38344 ;
  assign n38346 = n38345 ^ n37476 ;
  assign n38347 = n38346 ^ n36288 ;
  assign n38348 = n38347 ^ n38314 ;
  assign n38349 = n38348 ^ n38346 ;
  assign n38350 = ~n38339 & n38349 ;
  assign n38351 = n38350 ^ n38347 ;
  assign n38352 = n38351 ^ n36167 ;
  assign n38353 = n38352 ^ x438 ;
  assign n38357 = n38356 ^ n38353 ;
  assign n38338 = n38310 & n38332 ;
  assign n38358 = n38357 ^ n38338 ;
  assign n38309 = n38308 ^ n37926 ;
  assign n38335 = n38309 & n38334 ;
  assign n38336 = n38335 ^ n37926 ;
  assign n38337 = n38336 ^ n37922 ;
  assign n38389 = n38358 ^ n38337 ;
  assign n38848 = ~n37514 & ~n38389 ;
  assign n38849 = n38848 ^ n37922 ;
  assign n38850 = n38849 ^ n36855 ;
  assign n38851 = n38850 ^ n38819 ;
  assign n38852 = n38851 ^ n38849 ;
  assign n38853 = n38847 & ~n38852 ;
  assign n38854 = n38853 ^ n38850 ;
  assign n39028 = n38854 ^ n36816 ;
  assign n39224 = n39028 ^ x129 ;
  assign n39051 = n39050 ^ n39048 ;
  assign n39053 = ~n39051 & n39052 ;
  assign n39054 = n39053 ^ x130 ;
  assign n39225 = n39224 ^ n39054 ;
  assign n39226 = n39223 & n39225 ;
  assign n39055 = n39054 ^ n39028 ;
  assign n39056 = n39054 ^ x129 ;
  assign n39057 = ~n39055 & n39056 ;
  assign n39058 = n39057 ^ x129 ;
  assign n38384 = n38338 & n38357 ;
  assign n38378 = n38346 ^ n36167 ;
  assign n38379 = ~n38351 & n38378 ;
  assign n38380 = n38379 ^ n36167 ;
  assign n38373 = n37793 ^ n37791 ;
  assign n38367 = n38342 ^ n37791 ;
  assign n38370 = n38342 ^ n37476 ;
  assign n38371 = n38367 & n38370 ;
  assign n38368 = n37476 ^ n37472 ;
  assign n38372 = n38371 ^ n38368 ;
  assign n38374 = n38373 ^ n38372 ;
  assign n38375 = ~n36992 & n38374 ;
  assign n38376 = n38375 ^ n37472 ;
  assign n38377 = n38376 ^ n36162 ;
  assign n38381 = n38380 ^ n38377 ;
  assign n38382 = n38381 ^ x437 ;
  assign n38363 = n38356 ^ n38352 ;
  assign n38364 = n38356 ^ x438 ;
  assign n38365 = ~n38363 & n38364 ;
  assign n38366 = n38365 ^ x438 ;
  assign n38383 = n38382 ^ n38366 ;
  assign n38385 = n38384 ^ n38383 ;
  assign n38359 = n38358 ^ n38336 ;
  assign n38360 = n38337 & n38359 ;
  assign n38361 = n38360 ^ n37922 ;
  assign n38362 = n38361 ^ n37918 ;
  assign n38386 = n38385 ^ n38362 ;
  assign n38814 = n37510 & n38386 ;
  assign n38815 = n38814 ^ n37918 ;
  assign n38856 = n38815 ^ n36816 ;
  assign n38855 = n38849 ^ n38815 ;
  assign n38857 = n38856 ^ n38855 ;
  assign n38858 = n38854 & ~n38857 ;
  assign n38859 = n38858 ^ n38856 ;
  assign n39026 = n38859 ^ n36812 ;
  assign n39027 = n39026 ^ x128 ;
  assign n39227 = n39058 ^ n39027 ;
  assign n39228 = ~n39226 & n39227 ;
  assign n39059 = n39058 ^ n39026 ;
  assign n39060 = ~n39027 & n39059 ;
  assign n39061 = n39060 ^ x128 ;
  assign n39229 = n39061 ^ x143 ;
  assign n38816 = n38815 ^ n36812 ;
  assign n38860 = n38816 & ~n38859 ;
  assign n38861 = n38860 ^ n36812 ;
  assign n39023 = n38861 ^ n36867 ;
  assign n38691 = n38385 ^ n38361 ;
  assign n38470 = n38380 ^ n38376 ;
  assign n38471 = n38380 ^ n36162 ;
  assign n38472 = ~n38470 & n38471 ;
  assign n38473 = n38472 ^ n36162 ;
  assign n38405 = n38373 ^ n37472 ;
  assign n38406 = n38372 & n38405 ;
  assign n38407 = n38406 ^ n37472 ;
  assign n38403 = n37796 ^ n37794 ;
  assign n38404 = n38403 ^ n37469 ;
  assign n38466 = n38407 ^ n38404 ;
  assign n38467 = ~n36989 & ~n38466 ;
  assign n38468 = n38467 ^ n37469 ;
  assign n38469 = n38468 ^ n36303 ;
  assign n38565 = n38473 ^ n38469 ;
  assign n38641 = n38565 ^ x436 ;
  assign n38566 = n38381 ^ n38366 ;
  assign n38567 = n38382 & ~n38566 ;
  assign n38568 = n38567 ^ x437 ;
  assign n38642 = n38641 ^ n38568 ;
  assign n38640 = n38383 & n38384 ;
  assign n38689 = n38642 ^ n38640 ;
  assign n38692 = n38689 ^ n37918 ;
  assign n38693 = n38692 ^ n38689 ;
  assign n38694 = n38693 ^ n38361 ;
  assign n38695 = n38691 & ~n38694 ;
  assign n38696 = n38695 ^ n38692 ;
  assign n38862 = n38696 ^ n37913 ;
  assign n38863 = n37567 & ~n38862 ;
  assign n38864 = n38863 ^ n37913 ;
  assign n39024 = n39023 ^ n38864 ;
  assign n39230 = n39229 ^ n39024 ;
  assign n39231 = ~n39228 & ~n39230 ;
  assign n39025 = n39024 ^ x143 ;
  assign n39062 = n39061 ^ n39024 ;
  assign n39063 = ~n39025 & n39062 ;
  assign n39064 = n39063 ^ x143 ;
  assign n39232 = n39064 ^ x142 ;
  assign n38865 = n38864 ^ n38861 ;
  assign n38690 = n38689 ^ n37913 ;
  assign n38697 = n38690 & n38696 ;
  assign n38698 = n38697 ^ n37913 ;
  assign n38569 = n38568 ^ n38565 ;
  assign n38570 = n38568 ^ x436 ;
  assign n38571 = ~n38569 & n38570 ;
  assign n38572 = n38571 ^ x436 ;
  assign n38644 = n38572 ^ x435 ;
  assign n38408 = n38407 ^ n38403 ;
  assign n38409 = ~n38404 & ~n38408 ;
  assign n38410 = n38409 ^ n37469 ;
  assign n38401 = n37798 ^ n37797 ;
  assign n38402 = n38401 ^ n37614 ;
  assign n38463 = n38410 ^ n38402 ;
  assign n38464 = ~n36986 & n38463 ;
  assign n38465 = n38464 ^ n37614 ;
  assign n38562 = n38465 ^ n36158 ;
  assign n38474 = n38473 ^ n38468 ;
  assign n38475 = n38469 & n38474 ;
  assign n38476 = n38475 ^ n36303 ;
  assign n38563 = n38562 ^ n38476 ;
  assign n38645 = n38644 ^ n38563 ;
  assign n38643 = ~n38640 & ~n38642 ;
  assign n38687 = n38645 ^ n38643 ;
  assign n38688 = n38687 ^ n37909 ;
  assign n38866 = n38698 ^ n38688 ;
  assign n38867 = ~n37505 & n38866 ;
  assign n38868 = n38867 ^ n37909 ;
  assign n38869 = n38868 ^ n36867 ;
  assign n38870 = n38869 ^ n38861 ;
  assign n38871 = n38870 ^ n38868 ;
  assign n38872 = n38865 & ~n38871 ;
  assign n38873 = n38872 ^ n38869 ;
  assign n39021 = n38873 ^ n36734 ;
  assign n39233 = n39232 ^ n39021 ;
  assign n39234 = ~n39231 & n39233 ;
  assign n39022 = n39021 ^ x142 ;
  assign n39065 = n39064 ^ n39021 ;
  assign n39066 = ~n39022 & n39065 ;
  assign n39067 = n39066 ^ x142 ;
  assign n38699 = n38698 ^ n38687 ;
  assign n38700 = n38688 & ~n38699 ;
  assign n38701 = n38700 ^ n37909 ;
  assign n38809 = n38701 ^ n38006 ;
  assign n38411 = n38410 ^ n37614 ;
  assign n38412 = ~n38402 & ~n38411 ;
  assign n38413 = n38412 ^ n38401 ;
  assign n38399 = n37801 ^ n37799 ;
  assign n38400 = n38399 ^ n37465 ;
  assign n38481 = n38413 ^ n38400 ;
  assign n38482 = ~n36983 & ~n38481 ;
  assign n38483 = n38482 ^ n37465 ;
  assign n38560 = n38483 ^ n36154 ;
  assign n38477 = n38476 ^ n38465 ;
  assign n38478 = n38476 ^ n36158 ;
  assign n38479 = ~n38477 & ~n38478 ;
  assign n38480 = n38479 ^ n36158 ;
  assign n38561 = n38560 ^ n38480 ;
  assign n38647 = n38561 ^ x434 ;
  assign n38564 = n38563 ^ x435 ;
  assign n38573 = n38572 ^ n38563 ;
  assign n38574 = n38564 & ~n38573 ;
  assign n38575 = n38574 ^ x435 ;
  assign n38648 = n38647 ^ n38575 ;
  assign n38646 = ~n38643 & n38645 ;
  assign n38685 = n38648 ^ n38646 ;
  assign n38810 = n38809 ^ n38685 ;
  assign n38811 = n37500 & ~n38810 ;
  assign n38812 = n38811 ^ n38006 ;
  assign n38875 = n38812 ^ n36734 ;
  assign n38874 = n38868 ^ n38812 ;
  assign n38876 = n38875 ^ n38874 ;
  assign n38877 = ~n38873 & ~n38876 ;
  assign n38878 = n38877 ^ n38875 ;
  assign n39019 = n38878 ^ n36805 ;
  assign n39020 = n39019 ^ x141 ;
  assign n39235 = n39067 ^ n39020 ;
  assign n39236 = n39234 & ~n39235 ;
  assign n38813 = n38812 ^ n36805 ;
  assign n38879 = ~n38813 & ~n38878 ;
  assign n38880 = n38879 ^ n36805 ;
  assign n38686 = n38685 ^ n38006 ;
  assign n38702 = n38701 ^ n38685 ;
  assign n38703 = ~n38686 & ~n38702 ;
  assign n38704 = n38703 ^ n38006 ;
  assign n38804 = n38704 ^ n38097 ;
  assign n38576 = n38575 ^ n38561 ;
  assign n38577 = n38575 ^ x434 ;
  assign n38578 = n38576 & n38577 ;
  assign n38579 = n38578 ^ x434 ;
  assign n38484 = n38483 ^ n38480 ;
  assign n38416 = n37625 ^ n37465 ;
  assign n38414 = n38413 ^ n38399 ;
  assign n38415 = ~n38400 & ~n38414 ;
  assign n38417 = n38416 ^ n38415 ;
  assign n38397 = n37804 ^ n37802 ;
  assign n38459 = n38417 ^ n38397 ;
  assign n38460 = n36804 & ~n38459 ;
  assign n38461 = n38460 ^ n37625 ;
  assign n38485 = n38461 ^ n36154 ;
  assign n38486 = n38485 ^ n38461 ;
  assign n38487 = n38486 ^ n38480 ;
  assign n38488 = n38484 & n38487 ;
  assign n38489 = n38488 ^ n38485 ;
  assign n38558 = n38489 ^ n36150 ;
  assign n38559 = n38558 ^ x433 ;
  assign n38650 = n38579 ^ n38559 ;
  assign n38649 = n38646 & ~n38648 ;
  assign n38683 = n38650 ^ n38649 ;
  assign n38805 = n38804 ^ n38683 ;
  assign n38806 = n37496 & ~n38805 ;
  assign n38807 = n38806 ^ n38097 ;
  assign n38808 = n38807 ^ n36886 ;
  assign n39071 = n38880 ^ n38808 ;
  assign n39068 = n39067 ^ n39019 ;
  assign n39069 = n39020 & ~n39068 ;
  assign n39070 = n39069 ^ x141 ;
  assign n39072 = n39071 ^ n39070 ;
  assign n39237 = n39072 ^ x140 ;
  assign n39238 = n39236 & n39237 ;
  assign n38881 = n38880 ^ n38807 ;
  assign n38882 = ~n38808 & n38881 ;
  assign n38883 = n38882 ^ n36886 ;
  assign n39073 = n38883 ^ n36955 ;
  assign n38684 = n38683 ^ n38097 ;
  assign n38705 = n38704 ^ n38683 ;
  assign n38706 = n38684 & ~n38705 ;
  assign n38707 = n38706 ^ n38097 ;
  assign n38580 = n38579 ^ n38558 ;
  assign n38581 = n38559 & ~n38580 ;
  assign n38582 = n38581 ^ x433 ;
  assign n38652 = n38582 ^ x432 ;
  assign n38398 = n38397 ^ n37625 ;
  assign n38418 = n38398 & ~n38417 ;
  assign n38419 = n38418 ^ n38397 ;
  assign n38395 = n37807 ^ n37805 ;
  assign n38396 = n38395 ^ n37461 ;
  assign n38492 = n38419 ^ n38396 ;
  assign n38493 = ~n37072 & n38492 ;
  assign n38494 = n38493 ^ n37461 ;
  assign n38556 = n38494 ^ n36325 ;
  assign n38462 = n38461 ^ n36150 ;
  assign n38490 = n38462 & n38489 ;
  assign n38491 = n38490 ^ n36150 ;
  assign n38557 = n38556 ^ n38491 ;
  assign n38653 = n38652 ^ n38557 ;
  assign n38651 = n38649 & n38650 ;
  assign n38681 = n38653 ^ n38651 ;
  assign n38682 = n38681 ^ n38173 ;
  assign n38884 = n38707 ^ n38682 ;
  assign n38885 = ~n37491 & ~n38884 ;
  assign n38886 = n38885 ^ n38173 ;
  assign n39074 = n39073 ^ n38886 ;
  assign n39075 = n39074 ^ x140 ;
  assign n39076 = n39075 ^ n39070 ;
  assign n39077 = n39076 ^ n39074 ;
  assign n39078 = n39072 & n39077 ;
  assign n39079 = n39078 ^ n39075 ;
  assign n39239 = n39079 ^ x139 ;
  assign n39240 = n39238 & n39239 ;
  assign n38887 = n38886 ^ n38883 ;
  assign n38708 = n38707 ^ n38681 ;
  assign n38709 = n38682 & n38708 ;
  assign n38710 = n38709 ^ n38173 ;
  assign n38799 = n38710 ^ n38226 ;
  assign n38583 = n38582 ^ n38557 ;
  assign n38495 = n38494 ^ n38491 ;
  assign n38420 = n38419 ^ n38395 ;
  assign n38421 = ~n38396 & ~n38420 ;
  assign n38422 = n38421 ^ n37461 ;
  assign n38393 = n37809 ^ n37808 ;
  assign n38394 = n38393 ^ n37637 ;
  assign n38423 = n38422 ^ n38394 ;
  assign n38456 = ~n37068 & n38423 ;
  assign n38457 = n38456 ^ n37637 ;
  assign n38496 = n38457 ^ n36325 ;
  assign n38497 = n38496 ^ n38491 ;
  assign n38498 = n38497 ^ n38457 ;
  assign n38499 = n38495 & ~n38498 ;
  assign n38500 = n38499 ^ n38496 ;
  assign n38554 = n38500 ^ n36334 ;
  assign n38584 = n38554 ^ x432 ;
  assign n38585 = n38584 ^ n38557 ;
  assign n38586 = n38585 ^ n38554 ;
  assign n38587 = n38583 & ~n38586 ;
  assign n38588 = n38587 ^ n38584 ;
  assign n38655 = n38588 ^ x447 ;
  assign n38654 = n38651 & ~n38653 ;
  assign n38679 = n38655 ^ n38654 ;
  assign n38800 = n38799 ^ n38679 ;
  assign n38801 = ~n37487 & n38800 ;
  assign n38802 = n38801 ^ n38226 ;
  assign n38888 = n38802 ^ n36955 ;
  assign n38889 = n38888 ^ n38802 ;
  assign n38890 = n38889 ^ n38883 ;
  assign n38891 = ~n38887 & ~n38890 ;
  assign n38892 = n38891 ^ n38888 ;
  assign n39080 = n38892 ^ n37009 ;
  assign n39082 = n39080 ^ x139 ;
  assign n39081 = n39080 ^ n39074 ;
  assign n39083 = n39082 ^ n39081 ;
  assign n39084 = n39079 & ~n39083 ;
  assign n39085 = n39084 ^ n39082 ;
  assign n39241 = n39085 ^ x138 ;
  assign n39242 = n39240 & n39241 ;
  assign n38803 = n38802 ^ n37009 ;
  assign n38893 = n38803 & ~n38892 ;
  assign n38894 = n38893 ^ n37009 ;
  assign n39086 = n38894 ^ n37003 ;
  assign n38680 = n38679 ^ n38226 ;
  assign n38711 = n38710 ^ n38679 ;
  assign n38712 = n38680 & n38711 ;
  assign n38713 = n38712 ^ n38226 ;
  assign n38432 = n37811 ^ n37810 ;
  assign n38503 = n38432 ^ n37457 ;
  assign n38428 = n38422 ^ n38393 ;
  assign n38429 = n38422 ^ n37637 ;
  assign n38430 = ~n38428 & n38429 ;
  assign n38431 = n38430 ^ n37637 ;
  assign n38504 = n38503 ^ n38431 ;
  assign n38505 = ~n37064 & n38504 ;
  assign n38506 = n38505 ^ n37457 ;
  assign n38592 = n38506 ^ n36347 ;
  assign n38458 = n38457 ^ n36334 ;
  assign n38501 = n38458 & ~n38500 ;
  assign n38502 = n38501 ^ n36334 ;
  assign n38593 = n38592 ^ n38502 ;
  assign n38555 = n38554 ^ x447 ;
  assign n38589 = n38555 & ~n38588 ;
  assign n38590 = n38589 ^ x447 ;
  assign n38591 = n38590 ^ x446 ;
  assign n38657 = n38593 ^ n38591 ;
  assign n38656 = n38654 & n38655 ;
  assign n38677 = n38657 ^ n38656 ;
  assign n38678 = n38677 ^ n38265 ;
  assign n38795 = n38713 ^ n38678 ;
  assign n38796 = ~n37483 & n38795 ;
  assign n38797 = n38796 ^ n38265 ;
  assign n39087 = n39086 ^ n38797 ;
  assign n39089 = n39087 ^ x138 ;
  assign n39088 = n39087 ^ n39080 ;
  assign n39090 = n39089 ^ n39088 ;
  assign n39091 = n39085 & ~n39090 ;
  assign n39092 = n39091 ^ n39089 ;
  assign n39243 = n39092 ^ x137 ;
  assign n39244 = n39242 & ~n39243 ;
  assign n38798 = n38797 ^ n37003 ;
  assign n38895 = n38894 ^ n38797 ;
  assign n38896 = ~n38798 & ~n38895 ;
  assign n38897 = n38896 ^ n37003 ;
  assign n39016 = n38897 ^ n37001 ;
  assign n38714 = n38713 ^ n38677 ;
  assign n38715 = ~n38678 & n38714 ;
  assign n38716 = n38715 ^ n38265 ;
  assign n38790 = n38716 ^ n38278 ;
  assign n38507 = n38506 ^ n38502 ;
  assign n38433 = n38432 ^ n38431 ;
  assign n38426 = n37814 ^ n37812 ;
  assign n38434 = n38426 ^ n37457 ;
  assign n38435 = n38434 ^ n38426 ;
  assign n38436 = n38435 ^ n38431 ;
  assign n38437 = n38433 & ~n38436 ;
  assign n38438 = n38437 ^ n38434 ;
  assign n38508 = n38438 ^ n37892 ;
  assign n38509 = n37060 & ~n38508 ;
  assign n38510 = n38509 ^ n37892 ;
  assign n38511 = n38510 ^ n36347 ;
  assign n38512 = n38511 ^ n38502 ;
  assign n38513 = n38512 ^ n38510 ;
  assign n38514 = n38507 & ~n38513 ;
  assign n38515 = n38514 ^ n38511 ;
  assign n38598 = n38515 ^ n36509 ;
  assign n38594 = n38593 ^ n38590 ;
  assign n38595 = n38591 & ~n38594 ;
  assign n38596 = n38595 ^ x446 ;
  assign n38597 = n38596 ^ x445 ;
  assign n38659 = n38598 ^ n38597 ;
  assign n38658 = ~n38656 & ~n38657 ;
  assign n38717 = n38659 ^ n38658 ;
  assign n38791 = n38790 ^ n38717 ;
  assign n38792 = n37479 & n38791 ;
  assign n38793 = n38792 ^ n38278 ;
  assign n39017 = n39016 ^ n38793 ;
  assign n39094 = n39017 ^ x137 ;
  assign n39093 = n39087 ^ n39017 ;
  assign n39095 = n39094 ^ n39093 ;
  assign n39096 = ~n39092 & n39095 ;
  assign n39097 = n39096 ^ n39094 ;
  assign n39245 = n39097 ^ x136 ;
  assign n39246 = ~n39244 & ~n39245 ;
  assign n39018 = n39017 ^ x136 ;
  assign n39098 = ~n39018 & n39097 ;
  assign n39099 = n39098 ^ x136 ;
  assign n39247 = n39099 ^ x151 ;
  assign n38794 = n38793 ^ n37001 ;
  assign n38898 = n38897 ^ n38793 ;
  assign n38899 = ~n38794 & n38898 ;
  assign n38900 = n38899 ^ n37001 ;
  assign n39100 = n38900 ^ n36998 ;
  assign n38718 = n38717 ^ n38716 ;
  assign n38425 = n37817 ^ n37815 ;
  assign n38451 = n38425 ^ n37989 ;
  assign n38427 = n38426 ^ n37892 ;
  assign n38439 = n38427 & ~n38438 ;
  assign n38440 = n38439 ^ n37892 ;
  assign n38452 = n38451 ^ n38440 ;
  assign n38453 = ~n37156 & n38452 ;
  assign n38454 = n38453 ^ n37989 ;
  assign n38517 = n38454 ^ n36509 ;
  assign n38516 = n38510 ^ n38454 ;
  assign n38518 = n38517 ^ n38516 ;
  assign n38519 = ~n38515 & n38518 ;
  assign n38520 = n38519 ^ n38517 ;
  assign n38553 = n38520 ^ n36591 ;
  assign n38661 = n38553 ^ x444 ;
  assign n38599 = n38598 ^ n38596 ;
  assign n38600 = n38597 & n38599 ;
  assign n38601 = n38600 ^ x445 ;
  assign n38662 = n38661 ^ n38601 ;
  assign n38660 = n38658 & n38659 ;
  assign n38719 = n38662 ^ n38660 ;
  assign n38720 = n38719 ^ n38278 ;
  assign n38721 = n38720 ^ n38716 ;
  assign n38722 = n38721 ^ n38719 ;
  assign n38723 = n38718 & n38722 ;
  assign n38724 = n38723 ^ n38720 ;
  assign n38901 = n38724 ^ n38323 ;
  assign n38902 = ~n37597 & n38901 ;
  assign n38903 = n38902 ^ n38323 ;
  assign n39101 = n39100 ^ n38903 ;
  assign n39248 = n39247 ^ n39101 ;
  assign n39249 = ~n39246 & n39248 ;
  assign n39102 = n39101 ^ n39099 ;
  assign n38904 = n38903 ^ n38900 ;
  assign n38441 = n38440 ^ n38425 ;
  assign n38442 = n37820 ^ n37818 ;
  assign n38443 = n38442 ^ n37989 ;
  assign n38444 = n38443 ^ n38425 ;
  assign n38445 = n38444 ^ n38442 ;
  assign n38446 = ~n38441 & ~n38445 ;
  assign n38447 = n38446 ^ n38443 ;
  assign n38448 = n38447 ^ n38079 ;
  assign n38449 = n37056 & n38448 ;
  assign n38450 = n38449 ^ n38079 ;
  assign n38606 = n38450 ^ n36609 ;
  assign n38455 = n38454 ^ n36591 ;
  assign n38521 = n38455 & n38520 ;
  assign n38522 = n38521 ^ n36591 ;
  assign n38607 = n38606 ^ n38522 ;
  assign n38664 = n38607 ^ x443 ;
  assign n38602 = n38601 ^ n38553 ;
  assign n38603 = n38601 ^ x444 ;
  assign n38604 = n38602 & n38603 ;
  assign n38605 = n38604 ^ x444 ;
  assign n38665 = n38664 ^ n38605 ;
  assign n38663 = n38660 & n38662 ;
  assign n38725 = n38665 ^ n38663 ;
  assign n38727 = n38725 ^ n38323 ;
  assign n38726 = n38725 ^ n38719 ;
  assign n38728 = n38727 ^ n38726 ;
  assign n38729 = n38724 & ~n38728 ;
  assign n38730 = n38729 ^ n38727 ;
  assign n38786 = n38730 ^ n38344 ;
  assign n38787 = ~n37476 & ~n38786 ;
  assign n38788 = n38787 ^ n38344 ;
  assign n38905 = n38788 ^ n36998 ;
  assign n38906 = n38905 ^ n38788 ;
  assign n38907 = n38906 ^ n38900 ;
  assign n38908 = n38904 & n38907 ;
  assign n38909 = n38908 ^ n38905 ;
  assign n39103 = n38909 ^ n36996 ;
  assign n39104 = n39103 ^ x151 ;
  assign n39105 = n39104 ^ n39099 ;
  assign n39106 = n39105 ^ n39103 ;
  assign n39107 = n39102 & n39106 ;
  assign n39108 = n39107 ^ n39104 ;
  assign n39250 = n39108 ^ x150 ;
  assign n39251 = n39249 & n39250 ;
  assign n38789 = n38788 ^ n36996 ;
  assign n38910 = ~n38789 & n38909 ;
  assign n38911 = n38910 ^ n36996 ;
  assign n39109 = n38911 ^ n36992 ;
  assign n38608 = n38607 ^ n38605 ;
  assign n38523 = n38522 ^ n38450 ;
  assign n38524 = n38522 ^ n36609 ;
  assign n38525 = n38523 & n38524 ;
  assign n38526 = n38525 ^ n36609 ;
  assign n38609 = n38526 ^ n36634 ;
  assign n38527 = n37823 ^ n37821 ;
  assign n38529 = n38527 ^ n38079 ;
  assign n38528 = n38527 ^ n38442 ;
  assign n38530 = n38529 ^ n38528 ;
  assign n38531 = n38447 & n38530 ;
  assign n38532 = n38531 ^ n38529 ;
  assign n38533 = n38532 ^ n38155 ;
  assign n38534 = ~n37051 & ~n38533 ;
  assign n38535 = n38534 ^ n38155 ;
  assign n38610 = n38609 ^ n38535 ;
  assign n38611 = n38610 ^ x443 ;
  assign n38612 = n38611 ^ n38610 ;
  assign n38613 = n38612 ^ n38605 ;
  assign n38614 = n38608 & n38613 ;
  assign n38615 = n38614 ^ n38611 ;
  assign n38667 = n38615 ^ x442 ;
  assign n38666 = ~n38663 & ~n38665 ;
  assign n38675 = n38667 ^ n38666 ;
  assign n38732 = n38675 ^ n38344 ;
  assign n38731 = n38725 ^ n38675 ;
  assign n38733 = n38732 ^ n38731 ;
  assign n38734 = ~n38730 & n38733 ;
  assign n38735 = n38734 ^ n38732 ;
  assign n38782 = n38735 ^ n38374 ;
  assign n38783 = ~n37472 & ~n38782 ;
  assign n38784 = n38783 ^ n38374 ;
  assign n39110 = n39109 ^ n38784 ;
  assign n39112 = n39110 ^ x150 ;
  assign n39111 = n39110 ^ n39103 ;
  assign n39113 = n39112 ^ n39111 ;
  assign n39114 = n39108 & ~n39113 ;
  assign n39115 = n39114 ^ n39112 ;
  assign n39252 = n39115 ^ x149 ;
  assign n39253 = ~n39251 & ~n39252 ;
  assign n38785 = n38784 ^ n36992 ;
  assign n38912 = n38911 ^ n38784 ;
  assign n38913 = ~n38785 & ~n38912 ;
  assign n38914 = n38913 ^ n36992 ;
  assign n39116 = n38914 ^ n36989 ;
  assign n38676 = n38675 ^ n38374 ;
  assign n38736 = n38676 & n38735 ;
  assign n38737 = n38736 ^ n38374 ;
  assign n38777 = n38737 ^ n38466 ;
  assign n38536 = n38535 ^ n38526 ;
  assign n38542 = n37825 ^ n37824 ;
  assign n38538 = n38217 ^ n38155 ;
  assign n38537 = n38527 ^ n38217 ;
  assign n38539 = n38538 ^ n38537 ;
  assign n38540 = n38532 & n38539 ;
  assign n38541 = n38540 ^ n38538 ;
  assign n38543 = n38542 ^ n38541 ;
  assign n38544 = ~n37275 & ~n38543 ;
  assign n38545 = n38544 ^ n38217 ;
  assign n38546 = n38545 ^ n36634 ;
  assign n38547 = n38546 ^ n38545 ;
  assign n38548 = n38547 ^ n38526 ;
  assign n38549 = ~n38536 & ~n38548 ;
  assign n38550 = n38549 ^ n38546 ;
  assign n38551 = n38550 ^ n36650 ;
  assign n38617 = n38551 ^ x442 ;
  assign n38616 = n38610 ^ n38551 ;
  assign n38618 = n38617 ^ n38616 ;
  assign n38619 = n38615 & ~n38618 ;
  assign n38620 = n38619 ^ n38617 ;
  assign n38669 = n38620 ^ x441 ;
  assign n38668 = n38666 & ~n38667 ;
  assign n38673 = n38669 ^ n38668 ;
  assign n38778 = n38777 ^ n38673 ;
  assign n38779 = n37469 & ~n38778 ;
  assign n38780 = n38779 ^ n38466 ;
  assign n39117 = n39116 ^ n38780 ;
  assign n39119 = n39117 ^ x149 ;
  assign n39118 = n39117 ^ n39110 ;
  assign n39120 = n39119 ^ n39118 ;
  assign n39121 = n39115 & ~n39120 ;
  assign n39122 = n39121 ^ n39119 ;
  assign n39254 = n39122 ^ x148 ;
  assign n39255 = n39253 & ~n39254 ;
  assign n38781 = n38780 ^ n36989 ;
  assign n38915 = n38914 ^ n38780 ;
  assign n38916 = n38781 & ~n38915 ;
  assign n38917 = n38916 ^ n36989 ;
  assign n39123 = n38917 ^ n36986 ;
  assign n38674 = n38673 ^ n38466 ;
  assign n38738 = n38737 ^ n38673 ;
  assign n38739 = ~n38674 & ~n38738 ;
  assign n38740 = n38739 ^ n38466 ;
  assign n38772 = n38740 ^ n38463 ;
  assign n38670 = ~n38668 & ~n38669 ;
  assign n38633 = n37827 ^ n37826 ;
  assign n38634 = n38633 ^ n38250 ;
  assign n38635 = n38634 ^ n38542 ;
  assign n38631 = n38542 ^ n38217 ;
  assign n38632 = ~n38541 & ~n38631 ;
  assign n38636 = n38635 ^ n38632 ;
  assign n38637 = ~n37337 & n38636 ;
  assign n38626 = n38250 ^ n36689 ;
  assign n38627 = n38626 ^ n38545 ;
  assign n38623 = n36689 ^ n36650 ;
  assign n38624 = n38623 ^ n38250 ;
  assign n38628 = n38627 ^ n38624 ;
  assign n38629 = n38550 & ~n38628 ;
  assign n38622 = x441 ^ x440 ;
  assign n38625 = n38624 ^ n38622 ;
  assign n38630 = n38629 ^ n38625 ;
  assign n38638 = n38637 ^ n38630 ;
  assign n38552 = n38551 ^ x441 ;
  assign n38621 = n38552 & ~n38620 ;
  assign n38639 = n38638 ^ n38621 ;
  assign n38671 = n38670 ^ n38639 ;
  assign n38773 = n38772 ^ n38671 ;
  assign n38774 = n37614 & n38773 ;
  assign n38775 = n38774 ^ n38463 ;
  assign n39124 = n39123 ^ n38775 ;
  assign n39126 = n39124 ^ x148 ;
  assign n39125 = n39124 ^ n39117 ;
  assign n39127 = n39126 ^ n39125 ;
  assign n39128 = n39122 & ~n39127 ;
  assign n39129 = n39128 ^ n39126 ;
  assign n39256 = n39129 ^ x147 ;
  assign n39257 = ~n39255 & ~n39256 ;
  assign n38776 = n38775 ^ n36986 ;
  assign n38918 = n38917 ^ n38775 ;
  assign n38919 = ~n38776 & n38918 ;
  assign n38920 = n38919 ^ n36986 ;
  assign n39130 = n38920 ^ n36983 ;
  assign n38921 = n38481 ^ n38105 ;
  assign n38672 = n38671 ^ n38463 ;
  assign n38741 = n38740 ^ n38671 ;
  assign n38742 = ~n38672 & ~n38741 ;
  assign n38743 = n38742 ^ n38463 ;
  assign n38922 = n38921 ^ n38743 ;
  assign n38923 = n37465 & n38922 ;
  assign n38924 = n38923 ^ n38481 ;
  assign n39131 = n39130 ^ n38924 ;
  assign n39133 = n39131 ^ x147 ;
  assign n39132 = n39131 ^ n39124 ;
  assign n39134 = n39133 ^ n39132 ;
  assign n39135 = ~n39129 & n39134 ;
  assign n39136 = n39135 ^ n39133 ;
  assign n39258 = n39136 ^ x146 ;
  assign n39259 = ~n39257 & ~n39258 ;
  assign n38925 = n38924 ^ n38920 ;
  assign n38926 = n38924 ^ n36983 ;
  assign n38927 = ~n38925 & n38926 ;
  assign n38928 = n38927 ^ n36983 ;
  assign n39137 = n38928 ^ n36804 ;
  assign n38750 = n38106 ^ n38105 ;
  assign n38744 = n38743 ^ n38481 ;
  assign n38745 = n38459 ^ n38105 ;
  assign n38746 = n38745 ^ n38459 ;
  assign n38747 = n38746 ^ n38743 ;
  assign n38748 = n38744 & ~n38747 ;
  assign n38749 = n38748 ^ n38745 ;
  assign n38768 = n38750 ^ n38749 ;
  assign n38769 = n37625 & n38768 ;
  assign n38770 = n38769 ^ n38459 ;
  assign n39138 = n39137 ^ n38770 ;
  assign n39140 = n39138 ^ x146 ;
  assign n39139 = n39138 ^ n39131 ;
  assign n39141 = n39140 ^ n39139 ;
  assign n39142 = n39136 & ~n39141 ;
  assign n39143 = n39142 ^ n39140 ;
  assign n39260 = n39143 ^ x145 ;
  assign n39261 = ~n39259 & ~n39260 ;
  assign n38755 = n38107 ^ n38104 ;
  assign n38753 = n38492 ^ n38459 ;
  assign n38751 = n38750 ^ n38459 ;
  assign n38752 = n38749 & ~n38751 ;
  assign n38754 = n38753 ^ n38752 ;
  assign n38933 = n38755 ^ n38754 ;
  assign n38934 = ~n37461 & n38933 ;
  assign n38935 = n38934 ^ n38492 ;
  assign n38771 = n38770 ^ n36804 ;
  assign n38929 = n38928 ^ n38770 ;
  assign n38930 = ~n38771 & ~n38929 ;
  assign n38931 = n38930 ^ n36804 ;
  assign n38932 = n38931 ^ n37072 ;
  assign n39014 = n38935 ^ n38932 ;
  assign n39145 = n39014 ^ x145 ;
  assign n39144 = n39138 ^ n39014 ;
  assign n39146 = n39145 ^ n39144 ;
  assign n39147 = ~n39143 & n39146 ;
  assign n39148 = n39147 ^ n39145 ;
  assign n39262 = n39148 ^ x144 ;
  assign n39263 = ~n39261 & ~n39262 ;
  assign n39015 = n39014 ^ x144 ;
  assign n39149 = ~n39015 & n39148 ;
  assign n39150 = n39149 ^ x144 ;
  assign n39264 = n39150 ^ x159 ;
  assign n38936 = n38935 ^ n38931 ;
  assign n38937 = ~n38932 & ~n38936 ;
  assign n38938 = n38937 ^ n37072 ;
  assign n39151 = n38938 ^ n37068 ;
  assign n38392 = n38109 ^ n38108 ;
  assign n38756 = n38755 ^ n38392 ;
  assign n38757 = n38756 ^ n38492 ;
  assign n38758 = n38757 ^ n38392 ;
  assign n38759 = n38754 & ~n38758 ;
  assign n38760 = n38759 ^ n38756 ;
  assign n38939 = n38760 ^ n38423 ;
  assign n38940 = ~n37637 & ~n38939 ;
  assign n38941 = n38940 ^ n38423 ;
  assign n39152 = n39151 ^ n38941 ;
  assign n39265 = n39264 ^ n39152 ;
  assign n39266 = ~n39263 & ~n39265 ;
  assign n39153 = n39152 ^ n39150 ;
  assign n38942 = n38941 ^ n38938 ;
  assign n38424 = n38423 ^ n38392 ;
  assign n38761 = n38424 & n38760 ;
  assign n38762 = n38761 ^ n38423 ;
  assign n38391 = n38111 ^ n38110 ;
  assign n38763 = n38762 ^ n38391 ;
  assign n38764 = n38763 ^ n38504 ;
  assign n38765 = n37457 & ~n38764 ;
  assign n38766 = n38765 ^ n38504 ;
  assign n38943 = n38766 ^ n37068 ;
  assign n38944 = n38943 ^ n38938 ;
  assign n38945 = n38944 ^ n38766 ;
  assign n38946 = n38942 & n38945 ;
  assign n38947 = n38946 ^ n38943 ;
  assign n39154 = n38947 ^ n37064 ;
  assign n39155 = n39154 ^ x159 ;
  assign n39156 = n39155 ^ n39150 ;
  assign n39157 = n39156 ^ n39154 ;
  assign n39158 = ~n39153 & n39157 ;
  assign n39159 = n39158 ^ n39155 ;
  assign n39267 = n39159 ^ x158 ;
  assign n39268 = n39266 & ~n39267 ;
  assign n38767 = n38766 ^ n37064 ;
  assign n38948 = ~n38767 & n38947 ;
  assign n38949 = n38948 ^ n37064 ;
  assign n39160 = n38949 ^ n37060 ;
  assign n38955 = n38114 ^ n38112 ;
  assign n38951 = n38508 ^ n38504 ;
  assign n38950 = n38762 ^ n38508 ;
  assign n38952 = n38951 ^ n38950 ;
  assign n38953 = n38763 & n38952 ;
  assign n38954 = n38953 ^ n38951 ;
  assign n38956 = n38955 ^ n38954 ;
  assign n38957 = n37892 & ~n38956 ;
  assign n38958 = n38957 ^ n38508 ;
  assign n39161 = n39160 ^ n38958 ;
  assign n39163 = n39161 ^ x158 ;
  assign n39162 = n39161 ^ n39154 ;
  assign n39164 = n39163 ^ n39162 ;
  assign n39165 = ~n39159 & n39164 ;
  assign n39166 = n39165 ^ n39163 ;
  assign n39214 = n39166 ^ x157 ;
  assign n39276 = n39268 ^ n39214 ;
  assign n39308 = n39277 ^ n39276 ;
  assign n39269 = ~n39214 & n39268 ;
  assign n38959 = n38958 ^ n38949 ;
  assign n38960 = n38958 ^ n37060 ;
  assign n38961 = ~n38959 & ~n38960 ;
  assign n38962 = n38961 ^ n37060 ;
  assign n39167 = n38962 ^ n37156 ;
  assign n38968 = n38116 ^ n38115 ;
  assign n38964 = n38508 ^ n38452 ;
  assign n38963 = n38955 ^ n38452 ;
  assign n38965 = n38964 ^ n38963 ;
  assign n38966 = ~n38954 & ~n38965 ;
  assign n38967 = n38966 ^ n38964 ;
  assign n38969 = n38968 ^ n38967 ;
  assign n38970 = ~n37989 & ~n38969 ;
  assign n38971 = n38970 ^ n38452 ;
  assign n39168 = n39167 ^ n38971 ;
  assign n39170 = n39168 ^ x157 ;
  assign n39169 = n39168 ^ n39161 ;
  assign n39171 = n39170 ^ n39169 ;
  assign n39172 = ~n39166 & n39171 ;
  assign n39173 = n39172 ^ n39170 ;
  assign n39213 = n39173 ^ x156 ;
  assign n39279 = n39269 ^ n39213 ;
  assign n39278 = n39276 & n39277 ;
  assign n39280 = n39279 ^ n39278 ;
  assign n39309 = n39280 ^ n38183 ;
  assign n39310 = n39308 & ~n39309 ;
  assign n39270 = ~n39213 & ~n39269 ;
  assign n38972 = n38971 ^ n38962 ;
  assign n38973 = n38971 ^ n37156 ;
  assign n38974 = ~n38972 & ~n38973 ;
  assign n38975 = n38974 ^ n37156 ;
  assign n39174 = n38975 ^ n37056 ;
  assign n38981 = n38119 ^ n38117 ;
  assign n38977 = n38452 ^ n38448 ;
  assign n38976 = n38968 ^ n38448 ;
  assign n38978 = n38977 ^ n38976 ;
  assign n38979 = ~n38967 & n38978 ;
  assign n38980 = n38979 ^ n38977 ;
  assign n38982 = n38981 ^ n38980 ;
  assign n38983 = n38079 & n38982 ;
  assign n38984 = n38983 ^ n38448 ;
  assign n39175 = n39174 ^ n38984 ;
  assign n39177 = n39175 ^ x156 ;
  assign n39176 = n39175 ^ n39168 ;
  assign n39178 = n39177 ^ n39176 ;
  assign n39179 = n39173 & ~n39178 ;
  assign n39180 = n39179 ^ n39177 ;
  assign n39212 = n39180 ^ x155 ;
  assign n39284 = n39270 ^ n39212 ;
  assign n39281 = n39278 ^ n38183 ;
  assign n39282 = ~n39280 & ~n39281 ;
  assign n39283 = n39282 ^ n38183 ;
  assign n39285 = n39284 ^ n39283 ;
  assign n39311 = n39285 ^ n38826 ;
  assign n39312 = n39310 & ~n39311 ;
  assign n39271 = n39212 & ~n39270 ;
  assign n38985 = n38984 ^ n38975 ;
  assign n38986 = n38984 ^ n37056 ;
  assign n38987 = n38985 & n38986 ;
  assign n38988 = n38987 ^ n37056 ;
  assign n39181 = n38988 ^ n37051 ;
  assign n38994 = n38122 ^ n38120 ;
  assign n38990 = n38533 ^ n38448 ;
  assign n38989 = n38981 ^ n38533 ;
  assign n38991 = n38990 ^ n38989 ;
  assign n38992 = n38980 & n38991 ;
  assign n38993 = n38992 ^ n38990 ;
  assign n38995 = n38994 ^ n38993 ;
  assign n38996 = ~n38155 & n38995 ;
  assign n38997 = n38996 ^ n38533 ;
  assign n39182 = n39181 ^ n38997 ;
  assign n39184 = n39182 ^ x155 ;
  assign n39183 = n39182 ^ n39175 ;
  assign n39185 = n39184 ^ n39183 ;
  assign n39186 = n39180 & ~n39185 ;
  assign n39187 = n39186 ^ n39184 ;
  assign n39211 = n39187 ^ x154 ;
  assign n39290 = n39271 ^ n39211 ;
  assign n39286 = n39283 ^ n38826 ;
  assign n39287 = n39285 & ~n39286 ;
  assign n39288 = n39287 ^ n38826 ;
  assign n39289 = n39288 ^ n38836 ;
  assign n39313 = n39290 ^ n39289 ;
  assign n39314 = n39312 & ~n39313 ;
  assign n39008 = n38125 ^ n38123 ;
  assign n39004 = n38543 ^ n38533 ;
  assign n39003 = n38994 ^ n38543 ;
  assign n39005 = n39004 ^ n39003 ;
  assign n39006 = ~n38993 & n39005 ;
  assign n39007 = n39006 ^ n39004 ;
  assign n39009 = n39008 ^ n39007 ;
  assign n39010 = ~n38217 & ~n39009 ;
  assign n39011 = n39010 ^ n38543 ;
  assign n38998 = n38997 ^ n38988 ;
  assign n38999 = n38997 ^ n37051 ;
  assign n39000 = n38998 & n38999 ;
  assign n39001 = n39000 ^ n37051 ;
  assign n39002 = n39001 ^ n37275 ;
  assign n39012 = n39011 ^ n39002 ;
  assign n39189 = n39012 ^ x154 ;
  assign n39188 = n39182 ^ n39012 ;
  assign n39190 = n39189 ^ n39188 ;
  assign n39191 = ~n39187 & n39190 ;
  assign n39192 = n39191 ^ n39189 ;
  assign n39273 = n39192 ^ x153 ;
  assign n39272 = ~n39211 & n39271 ;
  assign n39295 = n39273 ^ n39272 ;
  assign n39291 = n39290 ^ n39288 ;
  assign n39292 = ~n39289 & ~n39291 ;
  assign n39293 = n39292 ^ n38836 ;
  assign n39294 = n39293 ^ n38821 ;
  assign n39315 = n39295 ^ n39294 ;
  assign n39316 = n39314 & ~n39315 ;
  assign n39296 = n39295 ^ n39293 ;
  assign n39297 = n39294 & ~n39296 ;
  assign n39298 = n39297 ^ n38821 ;
  assign n39317 = n39298 ^ n38817 ;
  assign n39274 = n39272 & n39273 ;
  assign n39204 = n38636 ^ n38126 ;
  assign n39205 = n39204 ^ n38128 ;
  assign n39206 = n39205 ^ n39008 ;
  assign n39202 = n39008 ^ n38543 ;
  assign n39203 = ~n39007 & n39202 ;
  assign n39207 = n39206 ^ n39203 ;
  assign n39208 = n38250 & n39207 ;
  assign n39198 = n37337 ^ n37275 ;
  assign n39199 = n39198 ^ n38636 ;
  assign n39197 = x153 ^ x152 ;
  assign n39200 = n39199 ^ n39197 ;
  assign n39194 = n39011 ^ n39001 ;
  assign n39195 = n39011 ^ n37275 ;
  assign n39196 = ~n39194 & n39195 ;
  assign n39201 = n39200 ^ n39196 ;
  assign n39209 = n39208 ^ n39201 ;
  assign n39013 = n39012 ^ x153 ;
  assign n39193 = ~n39013 & n39192 ;
  assign n39210 = n39209 ^ n39193 ;
  assign n39275 = n39274 ^ n39210 ;
  assign n39318 = n39317 ^ n39275 ;
  assign n39319 = n39316 & ~n39318 ;
  assign n39299 = n39298 ^ n39275 ;
  assign n39302 = n39275 ^ n38817 ;
  assign n39303 = n39299 & n39302 ;
  assign n39300 = n38817 ^ n38389 ;
  assign n39304 = n39303 ^ n39300 ;
  assign n38388 = n38136 ^ x135 ;
  assign n39320 = n39304 ^ n38388 ;
  assign n39321 = n39319 & n39320 ;
  assign n38390 = n38389 ^ n38388 ;
  assign n39305 = n38390 & n39304 ;
  assign n39306 = n39305 ^ n38389 ;
  assign n38387 = n38386 ^ n38189 ;
  assign n39307 = n39306 ^ n38387 ;
  assign n39322 = n39321 ^ n39307 ;
  assign n39323 = n39320 ^ n39319 ;
  assign n39324 = n39318 ^ n39316 ;
  assign n39325 = n39315 ^ n39314 ;
  assign n39326 = n39313 ^ n39312 ;
  assign n39327 = n39311 ^ n39310 ;
  assign n39328 = n39309 ^ n39308 ;
  assign n39373 = n39307 & n39321 ;
  assign n39344 = n39215 ^ n38189 ;
  assign n39340 = n38862 ^ n38386 ;
  assign n39338 = n39306 ^ n38189 ;
  assign n39339 = n38387 & n39338 ;
  assign n39341 = n39340 ^ n39339 ;
  assign n39374 = n39344 ^ n39341 ;
  assign n39375 = ~n39373 & n39374 ;
  assign n39348 = n39217 ^ n39216 ;
  assign n39342 = n38866 ^ n38862 ;
  assign n39343 = n39342 ^ n38866 ;
  assign n39345 = n39344 ^ n39343 ;
  assign n39346 = ~n39341 & n39345 ;
  assign n39347 = n39346 ^ n39342 ;
  assign n39376 = n39348 ^ n39347 ;
  assign n39377 = n39375 & n39376 ;
  assign n39336 = n39220 ^ n39218 ;
  assign n39350 = n39336 ^ n38866 ;
  assign n39349 = n39348 ^ n39336 ;
  assign n39351 = n39350 ^ n39349 ;
  assign n39352 = ~n39347 & ~n39351 ;
  assign n39353 = n39352 ^ n39350 ;
  assign n39378 = n39353 ^ n38810 ;
  assign n39379 = ~n39377 & ~n39378 ;
  assign n39357 = n39222 ^ n39221 ;
  assign n39337 = n39336 ^ n38810 ;
  assign n39354 = n39337 & n39353 ;
  assign n39335 = n38810 ^ n38805 ;
  assign n39355 = n39354 ^ n39335 ;
  assign n39380 = n39357 ^ n39355 ;
  assign n39381 = n39379 & n39380 ;
  assign n39333 = n39225 ^ n39223 ;
  assign n39356 = n39333 ^ n38805 ;
  assign n39358 = n39357 ^ n39356 ;
  assign n39359 = n39358 ^ n39333 ;
  assign n39360 = n39355 & n39359 ;
  assign n39361 = n39360 ^ n39356 ;
  assign n39382 = n39361 ^ n38884 ;
  assign n39383 = n39381 & n39382 ;
  assign n39364 = n39227 ^ n39226 ;
  assign n39334 = n39333 ^ n38884 ;
  assign n39362 = n39334 & ~n39361 ;
  assign n39332 = n38884 ^ n38800 ;
  assign n39363 = n39362 ^ n39332 ;
  assign n39384 = n39364 ^ n39363 ;
  assign n39385 = ~n39383 & n39384 ;
  assign n39368 = n39230 ^ n39228 ;
  assign n39365 = n39364 ^ n38800 ;
  assign n39366 = ~n39363 & ~n39365 ;
  assign n39331 = n38800 ^ n38795 ;
  assign n39367 = n39366 ^ n39331 ;
  assign n39386 = n39368 ^ n39367 ;
  assign n39387 = ~n39385 & n39386 ;
  assign n39369 = n39368 ^ n38795 ;
  assign n39370 = n39367 & ~n39369 ;
  assign n39330 = n38795 ^ n38791 ;
  assign n39371 = n39370 ^ n39330 ;
  assign n39329 = n39233 ^ n39231 ;
  assign n39372 = n39371 ^ n39329 ;
  assign n39388 = n39387 ^ n39372 ;
  assign n39389 = n39386 ^ n39385 ;
  assign n39390 = n39384 ^ n39383 ;
  assign n39391 = n39382 ^ n39381 ;
  assign n39392 = n39380 ^ n39379 ;
  assign n39393 = n39378 ^ n39377 ;
  assign n39394 = n39376 ^ n39375 ;
  assign n39395 = n39374 ^ n39373 ;
  assign n39438 = n39372 & n39387 ;
  assign n39402 = n39235 ^ n39234 ;
  assign n39439 = n39402 ^ n38901 ;
  assign n39403 = n39329 ^ n38791 ;
  assign n39404 = n39371 & ~n39403 ;
  assign n39405 = n39404 ^ n38791 ;
  assign n39440 = n39439 ^ n39405 ;
  assign n39441 = ~n39438 & ~n39440 ;
  assign n39406 = n39405 ^ n39402 ;
  assign n39400 = n39237 ^ n39236 ;
  assign n39407 = n39400 ^ n38901 ;
  assign n39408 = n39407 ^ n39402 ;
  assign n39409 = n39408 ^ n39400 ;
  assign n39410 = n39406 & ~n39409 ;
  assign n39411 = n39410 ^ n39407 ;
  assign n39442 = n39411 ^ n38786 ;
  assign n39443 = ~n39441 & n39442 ;
  assign n39414 = n39239 ^ n39238 ;
  assign n39401 = n39400 ^ n38786 ;
  assign n39412 = ~n39401 & ~n39411 ;
  assign n39399 = n38786 ^ n38782 ;
  assign n39413 = n39412 ^ n39399 ;
  assign n39444 = n39414 ^ n39413 ;
  assign n39445 = ~n39443 & n39444 ;
  assign n39418 = n39241 ^ n39240 ;
  assign n39415 = n39414 ^ n38782 ;
  assign n39416 = n39413 & ~n39415 ;
  assign n39398 = n38782 ^ n38778 ;
  assign n39417 = n39416 ^ n39398 ;
  assign n39446 = n39418 ^ n39417 ;
  assign n39447 = ~n39445 & ~n39446 ;
  assign n39422 = n39243 ^ n39242 ;
  assign n39419 = n39418 ^ n38778 ;
  assign n39420 = n39417 & ~n39419 ;
  assign n39397 = n38778 ^ n38773 ;
  assign n39421 = n39420 ^ n39397 ;
  assign n39448 = n39422 ^ n39421 ;
  assign n39449 = n39447 & ~n39448 ;
  assign n39427 = n39245 ^ n39244 ;
  assign n39425 = n38922 ^ n38773 ;
  assign n39423 = n39422 ^ n38773 ;
  assign n39424 = ~n39421 & ~n39423 ;
  assign n39426 = n39425 ^ n39424 ;
  assign n39450 = n39427 ^ n39426 ;
  assign n39451 = n39449 & n39450 ;
  assign n39396 = n39248 ^ n39246 ;
  assign n39452 = n39396 ^ n38768 ;
  assign n39428 = n39427 ^ n38922 ;
  assign n39429 = n39426 & ~n39428 ;
  assign n39430 = n39429 ^ n38922 ;
  assign n39453 = n39452 ^ n39430 ;
  assign n39454 = ~n39451 & ~n39453 ;
  assign n39435 = n39250 ^ n39249 ;
  assign n39436 = n39435 ^ n38933 ;
  assign n39431 = n39430 ^ n39396 ;
  assign n39432 = n39430 ^ n38768 ;
  assign n39433 = n39431 & n39432 ;
  assign n39434 = n39433 ^ n38768 ;
  assign n39437 = n39436 ^ n39434 ;
  assign n39455 = n39454 ^ n39437 ;
  assign n39456 = n39453 ^ n39451 ;
  assign n39457 = n39450 ^ n39449 ;
  assign n39458 = n39448 ^ n39447 ;
  assign n39459 = n39446 ^ n39445 ;
  assign n39460 = n39444 ^ n39443 ;
  assign n39461 = n39442 ^ n39441 ;
  assign n39462 = n39440 ^ n39438 ;
  assign n39514 = n39265 ^ n39263 ;
  assign n39515 = n39514 ^ n39009 ;
  assign n39507 = n39262 ^ n39261 ;
  assign n39508 = n39507 ^ n38995 ;
  assign n39464 = n39252 ^ n39251 ;
  assign n39465 = n39464 ^ n38939 ;
  assign n39466 = n39435 ^ n39434 ;
  assign n39467 = n39436 & ~n39466 ;
  assign n39468 = n39467 ^ n38933 ;
  assign n39471 = n39468 ^ n39464 ;
  assign n39475 = n39465 & n39471 ;
  assign n39472 = n38939 ^ n38764 ;
  assign n39476 = n39475 ^ n39472 ;
  assign n39481 = n38956 ^ n38764 ;
  assign n39477 = n39254 ^ n39253 ;
  assign n39480 = n39477 ^ n38956 ;
  assign n39482 = n39481 ^ n39480 ;
  assign n39483 = n39476 & ~n39482 ;
  assign n39484 = n39483 ^ n39481 ;
  assign n39489 = n38969 ^ n38956 ;
  assign n39485 = n39256 ^ n39255 ;
  assign n39488 = n39485 ^ n38969 ;
  assign n39490 = n39489 ^ n39488 ;
  assign n39491 = n39484 & ~n39490 ;
  assign n39492 = n39491 ^ n39489 ;
  assign n39496 = n39260 ^ n39259 ;
  assign n39498 = n39496 ^ n38969 ;
  assign n39493 = n39258 ^ n39257 ;
  assign n39497 = n39496 ^ n39493 ;
  assign n39499 = n39498 ^ n39497 ;
  assign n39500 = n39492 & n39499 ;
  assign n39501 = n39500 ^ n39498 ;
  assign n39504 = n39496 ^ n38982 ;
  assign n39505 = n39501 & n39504 ;
  assign n39506 = n39505 ^ n38982 ;
  assign n39511 = n39507 ^ n39506 ;
  assign n39512 = ~n39508 & n39511 ;
  assign n39513 = n39512 ^ n38995 ;
  assign n39521 = n39514 ^ n39513 ;
  assign n39522 = ~n39515 & n39521 ;
  assign n39518 = n39514 ^ n39266 ;
  assign n39519 = n39518 ^ n39267 ;
  assign n39520 = n39519 ^ n39207 ;
  assign n39523 = n39522 ^ n39520 ;
  assign n39463 = ~n39437 & ~n39454 ;
  assign n39469 = n39468 ^ n39465 ;
  assign n39470 = ~n39463 & n39469 ;
  assign n39478 = n39477 ^ n39476 ;
  assign n39479 = n39470 & n39478 ;
  assign n39486 = n39485 ^ n39484 ;
  assign n39487 = n39479 & n39486 ;
  assign n39494 = n39493 ^ n39492 ;
  assign n39495 = ~n39487 & n39494 ;
  assign n39502 = n39501 ^ n38982 ;
  assign n39503 = n39495 & n39502 ;
  assign n39509 = n39508 ^ n39506 ;
  assign n39510 = ~n39503 & ~n39509 ;
  assign n39516 = n39515 ^ n39513 ;
  assign n39517 = n39510 & ~n39516 ;
  assign n39524 = n39523 ^ n39517 ;
  assign n39525 = n39516 ^ n39510 ;
  assign n39526 = n39509 ^ n39503 ;
  assign n39527 = n39502 ^ n39495 ;
  assign n39528 = n39494 ^ n39487 ;
  assign n39529 = n39486 ^ n39479 ;
  assign n39530 = n39478 ^ n39470 ;
  assign n39531 = n39469 ^ n39463 ;
  assign n39541 = n37939 & ~n39308 ;
  assign n39542 = n39541 ^ n38131 ;
  assign n39580 = x359 & n39542 ;
  assign n39581 = n39580 ^ x358 ;
  assign n39543 = ~n37526 & ~n39542 ;
  assign n39582 = n39543 ^ n37531 ;
  assign n39544 = n37946 & n39309 ;
  assign n39545 = n39544 ^ n38183 ;
  assign n39583 = n39582 ^ n39545 ;
  assign n39584 = n39583 ^ n39580 ;
  assign n39585 = n39581 & ~n39584 ;
  assign n39586 = n39585 ^ x358 ;
  assign n39587 = n39586 ^ x357 ;
  assign n39546 = n39545 ^ n39543 ;
  assign n39547 = n39545 ^ n37531 ;
  assign n39548 = ~n39546 & n39547 ;
  assign n39549 = n39548 ^ n37531 ;
  assign n39588 = n39549 ^ n37523 ;
  assign n39538 = ~n37935 & n39311 ;
  assign n39539 = n39538 ^ n38826 ;
  assign n39589 = n39588 ^ n39539 ;
  assign n39590 = n39589 ^ n39586 ;
  assign n39591 = n39587 & n39590 ;
  assign n39592 = n39591 ^ x357 ;
  assign n39593 = n39592 ^ x356 ;
  assign n39540 = n39539 ^ n37523 ;
  assign n39550 = n39549 ^ n39539 ;
  assign n39551 = ~n39540 & n39550 ;
  assign n39552 = n39551 ^ n37523 ;
  assign n39594 = n39552 ^ n37518 ;
  assign n39553 = ~n37931 & n39313 ;
  assign n39554 = n39553 ^ n38836 ;
  assign n39595 = n39594 ^ n39554 ;
  assign n39596 = n39595 ^ n39592 ;
  assign n39597 = n39593 & ~n39596 ;
  assign n39598 = n39597 ^ x356 ;
  assign n39555 = n39554 ^ n39552 ;
  assign n39556 = n39554 ^ n37518 ;
  assign n39557 = ~n39555 & n39556 ;
  assign n39558 = n39557 ^ n37518 ;
  assign n39578 = n39558 ^ n37546 ;
  assign n39535 = ~n37957 & n39315 ;
  assign n39536 = n39535 ^ n38821 ;
  assign n39579 = n39578 ^ n39536 ;
  assign n39599 = n39598 ^ n39579 ;
  assign n39537 = n39536 ^ n37546 ;
  assign n39559 = n39558 ^ n39536 ;
  assign n39560 = n39537 & ~n39559 ;
  assign n39561 = n39560 ^ n37546 ;
  assign n39600 = n39561 ^ n37553 ;
  assign n39562 = ~n37926 & n39318 ;
  assign n39563 = n39562 ^ n38817 ;
  assign n39601 = n39600 ^ n39563 ;
  assign n39602 = n39601 ^ x355 ;
  assign n39603 = n39602 ^ n39598 ;
  assign n39604 = n39603 ^ n39601 ;
  assign n39605 = ~n39599 & n39604 ;
  assign n39606 = n39605 ^ n39602 ;
  assign n39731 = n39606 ^ x354 ;
  assign n39722 = n39542 ^ x359 ;
  assign n39723 = n39584 ^ x358 ;
  assign n39724 = n39722 & n39723 ;
  assign n39725 = n39590 ^ x357 ;
  assign n39726 = ~n39724 & n39725 ;
  assign n39727 = n39596 ^ x356 ;
  assign n39728 = ~n39726 & n39727 ;
  assign n39729 = n39599 ^ x355 ;
  assign n39730 = ~n39728 & ~n39729 ;
  assign n39762 = n39731 ^ n39730 ;
  assign n40152 = n39762 ^ n39372 ;
  assign n39763 = n39729 ^ n39728 ;
  assign n39764 = n39763 ^ n39386 ;
  assign n39766 = n39725 ^ n39724 ;
  assign n39767 = n39766 ^ n39382 ;
  assign n39768 = n39723 ^ n39722 ;
  assign n39769 = n39768 ^ n39380 ;
  assign n39564 = n39563 ^ n39561 ;
  assign n39565 = n39563 ^ n37553 ;
  assign n39566 = n39564 & ~n39565 ;
  assign n39567 = n39566 ^ n37553 ;
  assign n39575 = n39567 ^ n37514 ;
  assign n39532 = ~n37922 & ~n39320 ;
  assign n39533 = n39532 ^ n38389 ;
  assign n39576 = n39575 ^ n39533 ;
  assign n39577 = n39576 ^ x353 ;
  assign n39608 = n39576 ^ x354 ;
  assign n39607 = n39601 ^ n39576 ;
  assign n39609 = n39608 ^ n39607 ;
  assign n39610 = n39606 & ~n39609 ;
  assign n39611 = n39610 ^ n39608 ;
  assign n39612 = n39577 & ~n39611 ;
  assign n39613 = n39612 ^ x353 ;
  assign n39572 = n37918 & ~n39307 ;
  assign n39573 = n39572 ^ n38386 ;
  assign n39534 = n39533 ^ n37514 ;
  assign n39568 = n39567 ^ n39533 ;
  assign n39569 = n39534 & n39568 ;
  assign n39570 = n39569 ^ n37514 ;
  assign n39571 = n39570 ^ n37510 ;
  assign n39574 = n39573 ^ n39571 ;
  assign n39614 = n39613 ^ n39574 ;
  assign n39620 = ~n37913 & n39374 ;
  assign n39621 = n39620 ^ n38862 ;
  assign n39615 = n39573 ^ n39570 ;
  assign n39616 = n39573 ^ n37510 ;
  assign n39617 = n39615 & n39616 ;
  assign n39618 = n39617 ^ n37510 ;
  assign n39619 = n39618 ^ n37567 ;
  assign n39622 = n39621 ^ n39619 ;
  assign n39623 = n39622 ^ x352 ;
  assign n39624 = n39623 ^ n39613 ;
  assign n39625 = n39624 ^ n39622 ;
  assign n39626 = n39614 & n39625 ;
  assign n39627 = n39626 ^ n39623 ;
  assign n39633 = ~n37909 & n39376 ;
  assign n39634 = n39633 ^ n38866 ;
  assign n39628 = n39621 ^ n39618 ;
  assign n39629 = n39621 ^ n37567 ;
  assign n39630 = n39628 & ~n39629 ;
  assign n39631 = n39630 ^ n37567 ;
  assign n39632 = n39631 ^ n37505 ;
  assign n39635 = n39634 ^ n39632 ;
  assign n39637 = n39635 ^ x367 ;
  assign n39636 = n39635 ^ n39622 ;
  assign n39638 = n39637 ^ n39636 ;
  assign n39639 = n39627 & ~n39638 ;
  assign n39640 = n39639 ^ n39637 ;
  assign n39646 = n38006 & n39378 ;
  assign n39647 = n39646 ^ n38810 ;
  assign n39641 = n39634 ^ n39631 ;
  assign n39642 = n39634 ^ n37505 ;
  assign n39643 = ~n39641 & ~n39642 ;
  assign n39644 = n39643 ^ n37505 ;
  assign n39645 = n39644 ^ n37500 ;
  assign n39648 = n39647 ^ n39645 ;
  assign n39650 = n39648 ^ x366 ;
  assign n39649 = n39648 ^ n39635 ;
  assign n39651 = n39650 ^ n39649 ;
  assign n39652 = n39640 & ~n39651 ;
  assign n39653 = n39652 ^ n39650 ;
  assign n39659 = n38097 & ~n39380 ;
  assign n39660 = n39659 ^ n38805 ;
  assign n39654 = n39647 ^ n39644 ;
  assign n39655 = n39647 ^ n37500 ;
  assign n39656 = ~n39654 & ~n39655 ;
  assign n39657 = n39656 ^ n37500 ;
  assign n39658 = n39657 ^ n37496 ;
  assign n39661 = n39660 ^ n39658 ;
  assign n39663 = n39661 ^ x365 ;
  assign n39662 = n39661 ^ n39648 ;
  assign n39664 = n39663 ^ n39662 ;
  assign n39665 = ~n39653 & n39664 ;
  assign n39666 = n39665 ^ n39663 ;
  assign n39672 = ~n38173 & ~n39382 ;
  assign n39673 = n39672 ^ n38884 ;
  assign n39667 = n39660 ^ n39657 ;
  assign n39668 = n39660 ^ n37496 ;
  assign n39669 = n39667 & ~n39668 ;
  assign n39670 = n39669 ^ n37496 ;
  assign n39671 = n39670 ^ n37491 ;
  assign n39674 = n39673 ^ n39671 ;
  assign n39676 = n39674 ^ x364 ;
  assign n39675 = n39674 ^ n39661 ;
  assign n39677 = n39676 ^ n39675 ;
  assign n39678 = n39666 & ~n39677 ;
  assign n39679 = n39678 ^ n39676 ;
  assign n39685 = n38226 & n39384 ;
  assign n39686 = n39685 ^ n38800 ;
  assign n39680 = n39673 ^ n39670 ;
  assign n39681 = n39673 ^ n37491 ;
  assign n39682 = n39680 & n39681 ;
  assign n39683 = n39682 ^ n37491 ;
  assign n39684 = n39683 ^ n37487 ;
  assign n39687 = n39686 ^ n39684 ;
  assign n39689 = n39687 ^ x363 ;
  assign n39688 = n39687 ^ n39674 ;
  assign n39690 = n39689 ^ n39688 ;
  assign n39691 = ~n39679 & n39690 ;
  assign n39692 = n39691 ^ n39689 ;
  assign n39695 = n39686 ^ n39683 ;
  assign n39696 = n39686 ^ n37487 ;
  assign n39697 = n39695 & ~n39696 ;
  assign n39698 = n39697 ^ n37487 ;
  assign n39699 = n39698 ^ n37483 ;
  assign n39693 = n38265 & ~n39386 ;
  assign n39694 = n39693 ^ n38795 ;
  assign n39700 = n39699 ^ n39694 ;
  assign n39702 = n39700 ^ x362 ;
  assign n39701 = n39700 ^ n39687 ;
  assign n39703 = n39702 ^ n39701 ;
  assign n39704 = ~n39692 & n39703 ;
  assign n39705 = n39704 ^ n39702 ;
  assign n39711 = n38278 & ~n39372 ;
  assign n39712 = n39711 ^ n38791 ;
  assign n39706 = n39694 ^ n37483 ;
  assign n39707 = n39698 ^ n39694 ;
  assign n39708 = ~n39706 & n39707 ;
  assign n39709 = n39708 ^ n37483 ;
  assign n39710 = n39709 ^ n37479 ;
  assign n39713 = n39712 ^ n39710 ;
  assign n39715 = n39713 ^ x361 ;
  assign n39714 = n39713 ^ n39700 ;
  assign n39716 = n39715 ^ n39714 ;
  assign n39717 = ~n39705 & n39716 ;
  assign n39718 = n39717 ^ n39715 ;
  assign n39719 = n39718 ^ x360 ;
  assign n39720 = n39705 ^ x361 ;
  assign n39721 = n39692 ^ x362 ;
  assign n39732 = n39730 & n39731 ;
  assign n39733 = n39611 ^ x353 ;
  assign n39734 = ~n39732 & n39733 ;
  assign n39735 = n39614 ^ x352 ;
  assign n39736 = n39734 & ~n39735 ;
  assign n39737 = n39627 ^ x367 ;
  assign n39738 = n39736 & ~n39737 ;
  assign n39739 = n39640 ^ x366 ;
  assign n39740 = ~n39738 & n39739 ;
  assign n39741 = n39653 ^ x365 ;
  assign n39742 = ~n39740 & n39741 ;
  assign n39743 = n39666 ^ x364 ;
  assign n39744 = n39742 & ~n39743 ;
  assign n39745 = n39679 ^ x363 ;
  assign n39746 = ~n39744 & ~n39745 ;
  assign n39747 = ~n39721 & n39746 ;
  assign n39748 = ~n39720 & n39747 ;
  assign n39968 = n39719 & n39748 ;
  assign n39885 = n39713 ^ x360 ;
  assign n39886 = n39718 & ~n39885 ;
  assign n39887 = n39886 ^ x360 ;
  assign n39969 = n39887 ^ x375 ;
  assign n39797 = n39712 ^ n37479 ;
  assign n39798 = n39712 ^ n39709 ;
  assign n39799 = n39797 & n39798 ;
  assign n39800 = n39799 ^ n37479 ;
  assign n39883 = n39800 ^ n37597 ;
  assign n39801 = n38323 & ~n39440 ;
  assign n39802 = n39801 ^ n38901 ;
  assign n39884 = n39883 ^ n39802 ;
  assign n39970 = n39969 ^ n39884 ;
  assign n39971 = ~n39968 & ~n39970 ;
  assign n39888 = n39887 ^ n39884 ;
  assign n39803 = n39802 ^ n39800 ;
  assign n39794 = n38344 & ~n39442 ;
  assign n39795 = n39794 ^ n38786 ;
  assign n39804 = n39795 ^ n37597 ;
  assign n39805 = n39804 ^ n39795 ;
  assign n39806 = n39805 ^ n39800 ;
  assign n39807 = ~n39803 & ~n39806 ;
  assign n39808 = n39807 ^ n39804 ;
  assign n39889 = n39808 ^ n37476 ;
  assign n39890 = n39889 ^ x375 ;
  assign n39891 = n39890 ^ n39884 ;
  assign n39892 = n39891 ^ n39889 ;
  assign n39893 = n39888 & ~n39892 ;
  assign n39894 = n39893 ^ n39890 ;
  assign n39972 = n39894 ^ x374 ;
  assign n39973 = ~n39971 & n39972 ;
  assign n39796 = n39795 ^ n37476 ;
  assign n39809 = n39796 & ~n39808 ;
  assign n39810 = n39809 ^ n37476 ;
  assign n39895 = n39810 ^ n37472 ;
  assign n39791 = ~n38374 & n39444 ;
  assign n39792 = n39791 ^ n38782 ;
  assign n39896 = n39895 ^ n39792 ;
  assign n39898 = n39896 ^ x374 ;
  assign n39897 = n39896 ^ n39889 ;
  assign n39899 = n39898 ^ n39897 ;
  assign n39900 = n39894 & ~n39899 ;
  assign n39901 = n39900 ^ n39898 ;
  assign n39974 = n39901 ^ x373 ;
  assign n39975 = ~n39973 & ~n39974 ;
  assign n39793 = n39792 ^ n37472 ;
  assign n39811 = n39810 ^ n39792 ;
  assign n39812 = n39793 & ~n39811 ;
  assign n39813 = n39812 ^ n37472 ;
  assign n39880 = n39813 ^ n37469 ;
  assign n39788 = n38466 & n39446 ;
  assign n39789 = n39788 ^ n38778 ;
  assign n39881 = n39880 ^ n39789 ;
  assign n39903 = n39881 ^ x373 ;
  assign n39902 = n39896 ^ n39881 ;
  assign n39904 = n39903 ^ n39902 ;
  assign n39905 = n39901 & ~n39904 ;
  assign n39906 = n39905 ^ n39903 ;
  assign n39976 = n39906 ^ x372 ;
  assign n39977 = ~n39975 & ~n39976 ;
  assign n39790 = n39789 ^ n37469 ;
  assign n39814 = n39813 ^ n39789 ;
  assign n39815 = ~n39790 & ~n39814 ;
  assign n39816 = n39815 ^ n37469 ;
  assign n39878 = n39816 ^ n37614 ;
  assign n39785 = ~n38463 & n39448 ;
  assign n39786 = n39785 ^ n38773 ;
  assign n39879 = n39878 ^ n39786 ;
  assign n39978 = n39879 ^ x371 ;
  assign n39882 = n39881 ^ x372 ;
  assign n39907 = n39882 & ~n39906 ;
  assign n39908 = n39907 ^ x372 ;
  assign n39979 = n39978 ^ n39908 ;
  assign n39980 = n39977 & ~n39979 ;
  assign n39909 = n39908 ^ n39879 ;
  assign n39910 = n39908 ^ x371 ;
  assign n39911 = ~n39909 & n39910 ;
  assign n39912 = n39911 ^ x371 ;
  assign n39981 = n39912 ^ x370 ;
  assign n39787 = n39786 ^ n37614 ;
  assign n39817 = n39816 ^ n39786 ;
  assign n39818 = n39787 & ~n39817 ;
  assign n39819 = n39818 ^ n37614 ;
  assign n39913 = n39819 ^ n37465 ;
  assign n39820 = n38481 & ~n39450 ;
  assign n39821 = n39820 ^ n38922 ;
  assign n39914 = n39913 ^ n39821 ;
  assign n39982 = n39981 ^ n39914 ;
  assign n39983 = n39980 & ~n39982 ;
  assign n39915 = n39914 ^ n39912 ;
  assign n39822 = n39821 ^ n39819 ;
  assign n39782 = n38459 & ~n39453 ;
  assign n39783 = n39782 ^ n38768 ;
  assign n39823 = n39783 ^ n37465 ;
  assign n39824 = n39823 ^ n39783 ;
  assign n39825 = n39824 ^ n39819 ;
  assign n39826 = ~n39822 & n39825 ;
  assign n39827 = n39826 ^ n39823 ;
  assign n39876 = n39827 ^ n37625 ;
  assign n39916 = n39876 ^ x370 ;
  assign n39917 = n39916 ^ n39876 ;
  assign n39918 = n39917 ^ n39912 ;
  assign n39919 = ~n39915 & n39918 ;
  assign n39920 = n39919 ^ n39916 ;
  assign n39984 = n39920 ^ x369 ;
  assign n39985 = ~n39983 & n39984 ;
  assign n39877 = n39876 ^ x369 ;
  assign n39921 = n39877 & ~n39920 ;
  assign n39922 = n39921 ^ x369 ;
  assign n39784 = n39783 ^ n37625 ;
  assign n39828 = n39784 & ~n39827 ;
  assign n39829 = n39828 ^ n37625 ;
  assign n39779 = ~n38492 & n39437 ;
  assign n39780 = n39779 ^ n38933 ;
  assign n39781 = n39780 ^ n37461 ;
  assign n39874 = n39829 ^ n39781 ;
  assign n39875 = n39874 ^ x368 ;
  assign n39986 = n39922 ^ n39875 ;
  assign n39987 = n39985 & ~n39986 ;
  assign n39923 = n39922 ^ n39874 ;
  assign n39924 = ~n39875 & n39923 ;
  assign n39925 = n39924 ^ x368 ;
  assign n39988 = n39925 ^ x383 ;
  assign n39830 = n39829 ^ n39780 ;
  assign n39831 = ~n39781 & ~n39830 ;
  assign n39832 = n39831 ^ n37461 ;
  assign n39871 = n39832 ^ n37637 ;
  assign n39833 = ~n38423 & n39469 ;
  assign n39834 = n39833 ^ n38939 ;
  assign n39872 = n39871 ^ n39834 ;
  assign n39989 = n39988 ^ n39872 ;
  assign n39990 = ~n39987 & n39989 ;
  assign n39835 = n39834 ^ n39832 ;
  assign n39776 = ~n38504 & n39478 ;
  assign n39777 = n39776 ^ n38764 ;
  assign n39836 = n39777 ^ n37637 ;
  assign n39837 = n39836 ^ n39777 ;
  assign n39838 = n39837 ^ n39832 ;
  assign n39839 = ~n39835 & n39838 ;
  assign n39840 = n39839 ^ n39836 ;
  assign n39929 = n39840 ^ n37457 ;
  assign n39873 = n39872 ^ x383 ;
  assign n39926 = n39925 ^ n39872 ;
  assign n39927 = ~n39873 & n39926 ;
  assign n39928 = n39927 ^ x383 ;
  assign n39930 = n39929 ^ n39928 ;
  assign n39991 = n39930 ^ x382 ;
  assign n39992 = ~n39990 & n39991 ;
  assign n39931 = n39928 ^ x382 ;
  assign n39932 = ~n39930 & n39931 ;
  assign n39933 = n39932 ^ x382 ;
  assign n39778 = n39777 ^ n37457 ;
  assign n39841 = ~n39778 & ~n39840 ;
  assign n39842 = n39841 ^ n37457 ;
  assign n39773 = n38508 & n39486 ;
  assign n39774 = n39773 ^ n38956 ;
  assign n39775 = n39774 ^ n37892 ;
  assign n39869 = n39842 ^ n39775 ;
  assign n39870 = n39869 ^ x381 ;
  assign n39993 = n39933 ^ n39870 ;
  assign n39994 = ~n39992 & n39993 ;
  assign n39934 = n39933 ^ n39869 ;
  assign n39935 = ~n39870 & n39934 ;
  assign n39936 = n39935 ^ x381 ;
  assign n39995 = n39936 ^ x380 ;
  assign n39846 = ~n38452 & ~n39494 ;
  assign n39847 = n39846 ^ n38969 ;
  assign n39937 = n39847 ^ n37989 ;
  assign n39843 = n39842 ^ n39774 ;
  assign n39844 = ~n39775 & n39843 ;
  assign n39845 = n39844 ^ n37892 ;
  assign n39938 = n39937 ^ n39845 ;
  assign n39996 = n39995 ^ n39938 ;
  assign n39997 = n39994 & ~n39996 ;
  assign n39939 = n39938 ^ n39936 ;
  assign n39848 = n39847 ^ n39845 ;
  assign n39770 = ~n38448 & ~n39502 ;
  assign n39771 = n39770 ^ n38982 ;
  assign n39849 = n39771 ^ n37989 ;
  assign n39850 = n39849 ^ n39771 ;
  assign n39851 = n39850 ^ n39845 ;
  assign n39852 = n39848 & ~n39851 ;
  assign n39853 = n39852 ^ n39849 ;
  assign n39867 = n39853 ^ n38079 ;
  assign n39940 = n39867 ^ x380 ;
  assign n39941 = n39940 ^ n39867 ;
  assign n39942 = n39941 ^ n39936 ;
  assign n39943 = ~n39939 & n39942 ;
  assign n39944 = n39943 ^ n39940 ;
  assign n39998 = n39944 ^ x379 ;
  assign n39999 = n39997 & n39998 ;
  assign n39772 = n39771 ^ n38079 ;
  assign n39854 = n39772 & n39853 ;
  assign n39855 = n39854 ^ n38079 ;
  assign n39947 = n39855 ^ n38155 ;
  assign n39856 = n38533 & ~n39509 ;
  assign n39857 = n39856 ^ n38995 ;
  assign n39948 = n39947 ^ n39857 ;
  assign n40000 = n39948 ^ x378 ;
  assign n39868 = n39867 ^ x379 ;
  assign n39945 = ~n39868 & n39944 ;
  assign n39946 = n39945 ^ x379 ;
  assign n40001 = n40000 ^ n39946 ;
  assign n40002 = n39999 & n40001 ;
  assign n39949 = n39948 ^ n39946 ;
  assign n39863 = n38543 & ~n39516 ;
  assign n39864 = n39863 ^ n39009 ;
  assign n39858 = n39857 ^ n39855 ;
  assign n39859 = n39857 ^ n38155 ;
  assign n39860 = ~n39858 & ~n39859 ;
  assign n39861 = n39860 ^ n38155 ;
  assign n39862 = n39861 ^ n38217 ;
  assign n39865 = n39864 ^ n39862 ;
  assign n39950 = n39865 ^ x378 ;
  assign n39951 = n39950 ^ n39946 ;
  assign n39952 = n39951 ^ n39865 ;
  assign n39953 = n39949 & n39952 ;
  assign n39954 = n39953 ^ n39950 ;
  assign n39967 = n39954 ^ x377 ;
  assign n40005 = n40002 ^ n39967 ;
  assign n40006 = n40005 ^ n39374 ;
  assign n40040 = n40001 ^ n39999 ;
  assign n40007 = n39998 ^ n39997 ;
  assign n40008 = n40007 ^ n39320 ;
  assign n40009 = n39996 ^ n39994 ;
  assign n40010 = n40009 ^ n39318 ;
  assign n40029 = n39993 ^ n39992 ;
  assign n40011 = n39991 ^ n39990 ;
  assign n40012 = n40011 ^ n39313 ;
  assign n40013 = n39989 ^ n39987 ;
  assign n40014 = n40013 ^ n39311 ;
  assign n40016 = n39984 ^ n39983 ;
  assign n40017 = n39308 & ~n40016 ;
  assign n40015 = n39986 ^ n39985 ;
  assign n40018 = n40017 ^ n40015 ;
  assign n40019 = n40013 ^ n39309 ;
  assign n40020 = n40019 ^ n40013 ;
  assign n40021 = n40020 ^ n40015 ;
  assign n40022 = n40018 & n40021 ;
  assign n40023 = n40022 ^ n40019 ;
  assign n40024 = ~n40014 & n40023 ;
  assign n40025 = n40024 ^ n39311 ;
  assign n40026 = n40025 ^ n40011 ;
  assign n40027 = n40012 & ~n40026 ;
  assign n40028 = n40027 ^ n39313 ;
  assign n40030 = n40029 ^ n40028 ;
  assign n40031 = n40028 ^ n39315 ;
  assign n40032 = n40030 & n40031 ;
  assign n40033 = n40032 ^ n39315 ;
  assign n40034 = n40033 ^ n40009 ;
  assign n40035 = ~n40010 & n40034 ;
  assign n40036 = n40035 ^ n39318 ;
  assign n40037 = n40036 ^ n40007 ;
  assign n40038 = ~n40008 & ~n40037 ;
  assign n40039 = n40038 ^ n39320 ;
  assign n40041 = n40040 ^ n40039 ;
  assign n40042 = n40005 ^ n39307 ;
  assign n40043 = n40042 ^ n40005 ;
  assign n40044 = n40043 ^ n40039 ;
  assign n40045 = n40041 & n40044 ;
  assign n40046 = n40045 ^ n40042 ;
  assign n40047 = ~n40006 & ~n40046 ;
  assign n40048 = n40047 ^ n39374 ;
  assign n40003 = ~n39967 & ~n40002 ;
  assign n39964 = ~n38636 & ~n39523 ;
  assign n39960 = n38250 ^ n38217 ;
  assign n39961 = n39960 ^ n39207 ;
  assign n39959 = x377 ^ x376 ;
  assign n39962 = n39961 ^ n39959 ;
  assign n39956 = n39864 ^ n39861 ;
  assign n39957 = n39864 ^ n38217 ;
  assign n39958 = ~n39956 & n39957 ;
  assign n39963 = n39962 ^ n39958 ;
  assign n39965 = n39964 ^ n39963 ;
  assign n39866 = n39865 ^ x377 ;
  assign n39955 = ~n39866 & n39954 ;
  assign n39966 = n39965 ^ n39955 ;
  assign n40004 = n40003 ^ n39966 ;
  assign n40049 = n40048 ^ n40004 ;
  assign n40050 = n39722 ^ n39376 ;
  assign n40051 = n40050 ^ n39722 ;
  assign n40052 = n40051 ^ n40004 ;
  assign n40053 = n40049 & ~n40052 ;
  assign n40054 = n40053 ^ n40050 ;
  assign n40056 = n39380 ^ n39378 ;
  assign n40055 = n39722 ^ n39380 ;
  assign n40057 = n40056 ^ n40055 ;
  assign n40058 = ~n40054 & n40057 ;
  assign n40059 = n40058 ^ n40056 ;
  assign n40060 = n39769 & ~n40059 ;
  assign n40061 = n40060 ^ n39380 ;
  assign n40062 = n40061 ^ n39766 ;
  assign n40063 = n39767 & ~n40062 ;
  assign n40064 = n40063 ^ n39382 ;
  assign n39765 = n39727 ^ n39726 ;
  assign n40065 = n40064 ^ n39765 ;
  assign n40067 = n39386 ^ n39384 ;
  assign n40066 = n40064 ^ n39386 ;
  assign n40068 = n40067 ^ n40066 ;
  assign n40069 = n40065 & ~n40068 ;
  assign n40070 = n40069 ^ n40067 ;
  assign n40071 = ~n39764 & ~n40070 ;
  assign n40072 = n40071 ^ n39386 ;
  assign n40153 = n40152 ^ n40072 ;
  assign n40154 = ~n38791 & n40153 ;
  assign n40155 = n40154 ^ n39372 ;
  assign n40156 = n40155 ^ n38278 ;
  assign n40157 = n40070 ^ n39763 ;
  assign n40158 = ~n38795 & ~n40157 ;
  assign n40159 = n40158 ^ n39386 ;
  assign n40160 = n40159 ^ n38265 ;
  assign n40161 = n40065 ^ n39384 ;
  assign n40162 = ~n38800 & ~n40161 ;
  assign n40163 = n40162 ^ n39384 ;
  assign n40164 = n40163 ^ n38226 ;
  assign n40165 = n40061 ^ n39767 ;
  assign n40166 = n38884 & ~n40165 ;
  assign n40167 = n40166 ^ n39382 ;
  assign n40168 = n40167 ^ n38173 ;
  assign n40169 = n40059 ^ n39768 ;
  assign n40170 = n38805 & n40169 ;
  assign n40171 = n40170 ^ n39380 ;
  assign n40172 = n40171 ^ n38097 ;
  assign n40245 = n40054 ^ n39378 ;
  assign n40246 = n38810 & n40245 ;
  assign n40247 = n40246 ^ n39378 ;
  assign n40173 = n40048 ^ n39376 ;
  assign n40174 = n40173 ^ n40004 ;
  assign n40175 = ~n38866 & ~n40174 ;
  assign n40176 = n40175 ^ n39376 ;
  assign n40177 = n40176 ^ n37909 ;
  assign n40178 = n40046 ^ n39374 ;
  assign n40179 = n38862 & n40178 ;
  assign n40180 = n40179 ^ n39374 ;
  assign n40181 = n40180 ^ n37913 ;
  assign n40182 = n40040 ^ n39307 ;
  assign n40183 = n40182 ^ n40039 ;
  assign n40184 = ~n38386 & n40183 ;
  assign n40185 = n40184 ^ n39307 ;
  assign n40186 = n40185 ^ n37918 ;
  assign n40187 = n40036 ^ n40008 ;
  assign n40188 = n38389 & ~n40187 ;
  assign n40189 = n40188 ^ n39320 ;
  assign n40190 = n40189 ^ n37922 ;
  assign n40191 = n40030 ^ n39315 ;
  assign n40192 = ~n38821 & ~n40191 ;
  assign n40193 = n40192 ^ n39315 ;
  assign n40194 = n40193 ^ n37957 ;
  assign n40215 = n40025 ^ n40012 ;
  assign n40216 = ~n38836 & n40215 ;
  assign n40217 = n40216 ^ n39313 ;
  assign n40195 = n40016 ^ n39276 ;
  assign n40196 = n40195 ^ n39277 ;
  assign n40197 = n39277 & n40196 ;
  assign n40198 = n40197 ^ n39308 ;
  assign n40199 = n37939 & ~n40198 ;
  assign n40200 = n40199 ^ n37946 ;
  assign n40204 = n40199 ^ n39280 ;
  assign n40201 = n40015 ^ n39309 ;
  assign n40202 = n40201 ^ n40017 ;
  assign n40203 = ~n38183 & n40202 ;
  assign n40205 = n40204 ^ n40203 ;
  assign n40206 = n40200 & n40205 ;
  assign n40207 = n40206 ^ n37946 ;
  assign n40208 = n40207 ^ n37935 ;
  assign n40209 = n40023 ^ n39311 ;
  assign n40210 = n38826 & ~n40209 ;
  assign n40211 = n40210 ^ n39311 ;
  assign n40212 = n40211 ^ n40207 ;
  assign n40213 = ~n40208 & ~n40212 ;
  assign n40214 = n40213 ^ n37935 ;
  assign n40218 = n40217 ^ n40214 ;
  assign n40219 = n40217 ^ n37931 ;
  assign n40220 = n40218 & ~n40219 ;
  assign n40221 = n40220 ^ n37931 ;
  assign n40222 = n40221 ^ n40193 ;
  assign n40223 = ~n40194 & n40222 ;
  assign n40224 = n40223 ^ n37957 ;
  assign n40225 = n40224 ^ n37926 ;
  assign n40226 = n40033 ^ n39318 ;
  assign n40227 = n40226 ^ n40009 ;
  assign n40228 = n38817 & ~n40227 ;
  assign n40229 = n40228 ^ n39318 ;
  assign n40230 = n40229 ^ n40224 ;
  assign n40231 = n40225 & n40230 ;
  assign n40232 = n40231 ^ n37926 ;
  assign n40233 = n40232 ^ n40189 ;
  assign n40234 = n40190 & ~n40233 ;
  assign n40235 = n40234 ^ n37922 ;
  assign n40236 = n40235 ^ n40185 ;
  assign n40237 = ~n40186 & ~n40236 ;
  assign n40238 = n40237 ^ n37918 ;
  assign n40239 = n40238 ^ n40180 ;
  assign n40240 = ~n40181 & ~n40239 ;
  assign n40241 = n40240 ^ n37913 ;
  assign n40242 = n40241 ^ n40176 ;
  assign n40243 = ~n40177 & n40242 ;
  assign n40244 = n40243 ^ n37909 ;
  assign n40248 = n40247 ^ n40244 ;
  assign n40249 = n40171 ^ n38006 ;
  assign n40250 = n40249 ^ n40171 ;
  assign n40251 = n40250 ^ n40244 ;
  assign n40252 = n40248 & ~n40251 ;
  assign n40253 = n40252 ^ n40249 ;
  assign n40254 = ~n40172 & n40253 ;
  assign n40255 = n40254 ^ n38097 ;
  assign n40256 = n40255 ^ n40167 ;
  assign n40257 = n40168 & n40256 ;
  assign n40258 = n40257 ^ n38173 ;
  assign n40259 = n40258 ^ n40163 ;
  assign n40260 = n40164 & n40259 ;
  assign n40261 = n40260 ^ n38226 ;
  assign n40262 = n40261 ^ n40159 ;
  assign n40263 = ~n40160 & n40262 ;
  assign n40264 = n40263 ^ n38265 ;
  assign n40265 = n40264 ^ n40155 ;
  assign n40266 = ~n40156 & n40265 ;
  assign n40267 = n40266 ^ n38278 ;
  assign n40315 = n40267 ^ n38323 ;
  assign n40073 = n40072 ^ n39762 ;
  assign n40074 = n39440 ^ n39372 ;
  assign n40075 = n40074 ^ n39440 ;
  assign n40076 = n40075 ^ n39762 ;
  assign n40077 = n40073 & ~n40076 ;
  assign n40078 = n40077 ^ n40074 ;
  assign n39760 = n39733 ^ n39732 ;
  assign n40148 = n40078 ^ n39760 ;
  assign n40149 = ~n38901 & n40148 ;
  assign n40150 = n40149 ^ n39440 ;
  assign n40316 = n40315 ^ n40150 ;
  assign n40317 = n40316 ^ x87 ;
  assign n40318 = n40264 ^ n40156 ;
  assign n40319 = n40318 ^ x72 ;
  assign n40401 = n40261 ^ n40160 ;
  assign n40320 = n40258 ^ n38226 ;
  assign n40321 = n40320 ^ n40163 ;
  assign n40322 = n40321 ^ x74 ;
  assign n40378 = n40244 ^ n38006 ;
  assign n40379 = n40378 ^ n40247 ;
  assign n40323 = n40241 ^ n40177 ;
  assign n40324 = n40323 ^ x78 ;
  assign n40325 = n40238 ^ n37913 ;
  assign n40326 = n40325 ^ n40180 ;
  assign n40327 = n40326 ^ x79 ;
  assign n40365 = n40235 ^ n37918 ;
  assign n40366 = n40365 ^ n40185 ;
  assign n40328 = n40232 ^ n37922 ;
  assign n40329 = n40328 ^ n40189 ;
  assign n40330 = n40329 ^ x65 ;
  assign n40332 = n40214 ^ n37931 ;
  assign n40333 = n40332 ^ n40217 ;
  assign n40334 = n40333 ^ x68 ;
  assign n40343 = n40211 ^ n40208 ;
  assign n40336 = n39276 ^ n38130 ;
  assign n40337 = n40336 ^ n40197 ;
  assign n40338 = x71 & ~n40337 ;
  assign n40335 = n40205 ^ n37946 ;
  assign n40339 = n40338 ^ n40335 ;
  assign n40340 = n40338 ^ x70 ;
  assign n40341 = n40339 & n40340 ;
  assign n40342 = n40341 ^ x70 ;
  assign n40344 = n40343 ^ n40342 ;
  assign n40347 = n40342 ^ x69 ;
  assign n40348 = n40344 & n40347 ;
  assign n40345 = n40333 ^ x69 ;
  assign n40349 = n40348 ^ n40345 ;
  assign n40350 = n40334 & ~n40349 ;
  assign n40351 = n40350 ^ x68 ;
  assign n40352 = n40351 ^ x67 ;
  assign n40353 = n40221 ^ n37957 ;
  assign n40354 = n40353 ^ n40193 ;
  assign n40355 = n40354 ^ n40351 ;
  assign n40356 = n40352 & ~n40355 ;
  assign n40357 = n40356 ^ x67 ;
  assign n40331 = n40229 ^ n40225 ;
  assign n40358 = n40357 ^ n40331 ;
  assign n40359 = n40357 ^ x66 ;
  assign n40360 = ~n40358 & n40359 ;
  assign n40361 = n40360 ^ x66 ;
  assign n40362 = n40361 ^ n40329 ;
  assign n40363 = ~n40330 & n40362 ;
  assign n40364 = n40363 ^ x65 ;
  assign n40367 = n40366 ^ n40364 ;
  assign n40368 = n40326 ^ x64 ;
  assign n40369 = n40368 ^ n40326 ;
  assign n40370 = n40369 ^ n40364 ;
  assign n40371 = ~n40367 & n40370 ;
  assign n40372 = n40371 ^ n40368 ;
  assign n40373 = ~n40327 & n40372 ;
  assign n40374 = n40373 ^ x79 ;
  assign n40375 = n40374 ^ n40323 ;
  assign n40376 = n40324 & ~n40375 ;
  assign n40377 = n40376 ^ x78 ;
  assign n40380 = n40379 ^ n40377 ;
  assign n40381 = n40253 ^ n38097 ;
  assign n40382 = n40381 ^ x77 ;
  assign n40383 = n40382 ^ n40377 ;
  assign n40384 = n40383 ^ n40381 ;
  assign n40385 = n40380 & n40384 ;
  assign n40386 = n40385 ^ n40382 ;
  assign n40387 = n40255 ^ n38173 ;
  assign n40388 = n40387 ^ n40167 ;
  assign n40390 = n40388 ^ x76 ;
  assign n40389 = n40388 ^ n40381 ;
  assign n40391 = n40390 ^ n40389 ;
  assign n40392 = n40386 & ~n40391 ;
  assign n40393 = n40392 ^ n40390 ;
  assign n40395 = n40321 ^ x75 ;
  assign n40394 = n40388 ^ n40321 ;
  assign n40396 = n40395 ^ n40394 ;
  assign n40397 = ~n40393 & n40396 ;
  assign n40398 = n40397 ^ n40395 ;
  assign n40399 = ~n40322 & n40398 ;
  assign n40400 = n40399 ^ x74 ;
  assign n40402 = n40401 ^ n40400 ;
  assign n40403 = n40318 ^ x73 ;
  assign n40404 = n40403 ^ n40318 ;
  assign n40405 = n40404 ^ n40400 ;
  assign n40406 = n40402 & n40405 ;
  assign n40407 = n40406 ^ n40403 ;
  assign n40408 = ~n40319 & n40407 ;
  assign n40409 = n40408 ^ x72 ;
  assign n40410 = n40409 ^ n40316 ;
  assign n40411 = ~n40317 & n40410 ;
  assign n40412 = n40411 ^ x87 ;
  assign n40151 = n40150 ^ n38323 ;
  assign n40268 = n40267 ^ n40150 ;
  assign n40269 = ~n40151 & n40268 ;
  assign n40270 = n40269 ^ n38323 ;
  assign n39759 = n39735 ^ n39734 ;
  assign n40143 = n39759 ^ n39442 ;
  assign n39761 = n39760 ^ n39440 ;
  assign n40079 = ~n39761 & n40078 ;
  assign n40080 = n40079 ^ n39440 ;
  assign n40144 = n40143 ^ n40080 ;
  assign n40145 = n38786 & n40144 ;
  assign n40146 = n40145 ^ n39442 ;
  assign n40147 = n40146 ^ n38344 ;
  assign n40313 = n40270 ^ n40147 ;
  assign n40314 = n40313 ^ x86 ;
  assign n40532 = n40412 ^ n40314 ;
  assign n40491 = n40337 ^ x71 ;
  assign n40492 = n40335 ^ x70 ;
  assign n40493 = n40492 ^ n40338 ;
  assign n40494 = n40491 & n40493 ;
  assign n40495 = n40343 ^ x69 ;
  assign n40496 = n40495 ^ n40342 ;
  assign n40497 = ~n40494 & ~n40496 ;
  assign n40498 = n40349 ^ x68 ;
  assign n40499 = ~n40497 & ~n40498 ;
  assign n40500 = n40355 ^ x67 ;
  assign n40501 = n40499 & ~n40500 ;
  assign n40502 = n40331 ^ x66 ;
  assign n40503 = n40502 ^ n40357 ;
  assign n40504 = n40501 & ~n40503 ;
  assign n40505 = n40361 ^ x65 ;
  assign n40506 = n40505 ^ n40329 ;
  assign n40507 = ~n40504 & ~n40506 ;
  assign n40508 = n40366 ^ x64 ;
  assign n40509 = n40508 ^ n40364 ;
  assign n40510 = ~n40507 & ~n40509 ;
  assign n40511 = n40372 ^ x79 ;
  assign n40512 = ~n40510 & ~n40511 ;
  assign n40513 = n40374 ^ x78 ;
  assign n40514 = n40513 ^ n40323 ;
  assign n40515 = ~n40512 & ~n40514 ;
  assign n40516 = n40377 ^ x77 ;
  assign n40517 = n40516 ^ n40379 ;
  assign n40518 = ~n40515 & ~n40517 ;
  assign n40519 = n40386 ^ x76 ;
  assign n40520 = n40518 & ~n40519 ;
  assign n40521 = n40393 ^ x75 ;
  assign n40522 = ~n40520 & ~n40521 ;
  assign n40523 = n40398 ^ x74 ;
  assign n40524 = ~n40522 & ~n40523 ;
  assign n40525 = n40400 ^ x73 ;
  assign n40526 = n40525 ^ n40401 ;
  assign n40527 = ~n40524 & n40526 ;
  assign n40528 = n40407 ^ x72 ;
  assign n40529 = n40527 & n40528 ;
  assign n40530 = n40409 ^ n40317 ;
  assign n40531 = n40529 & n40530 ;
  assign n40569 = n40532 ^ n40531 ;
  assign n40688 = n40569 ^ n40196 ;
  assign n40689 = n39308 & ~n40688 ;
  assign n40690 = n40689 ^ n40195 ;
  assign n40900 = n40690 ^ x295 ;
  assign n40835 = x295 & n40690 ;
  assign n40901 = n40835 ^ x294 ;
  assign n40691 = n39277 & ~n40690 ;
  assign n40833 = n40691 ^ n38183 ;
  assign n40271 = n40270 ^ n40146 ;
  assign n40272 = ~n40147 & n40271 ;
  assign n40273 = n40272 ^ n38344 ;
  assign n40416 = n40273 ^ n38374 ;
  assign n40087 = n39737 ^ n39736 ;
  assign n40081 = n40080 ^ n39759 ;
  assign n40082 = n39444 ^ n39442 ;
  assign n40083 = n40082 ^ n39444 ;
  assign n40084 = n40083 ^ n39759 ;
  assign n40085 = n40081 & ~n40084 ;
  assign n40086 = n40085 ^ n40082 ;
  assign n40139 = n40087 ^ n40086 ;
  assign n40140 = n38782 & ~n40139 ;
  assign n40141 = n40140 ^ n39444 ;
  assign n40417 = n40416 ^ n40141 ;
  assign n40534 = n40417 ^ x85 ;
  assign n40413 = n40412 ^ n40313 ;
  assign n40414 = ~n40314 & n40413 ;
  assign n40415 = n40414 ^ x86 ;
  assign n40535 = n40534 ^ n40415 ;
  assign n40533 = n40531 & n40532 ;
  assign n40572 = n40535 ^ n40533 ;
  assign n40570 = ~n40196 & ~n40569 ;
  assign n40571 = n40570 ^ n40202 ;
  assign n40692 = n40572 ^ n40571 ;
  assign n40693 = ~n39309 & n40692 ;
  assign n40694 = n40693 ^ n40202 ;
  assign n40834 = n40833 ^ n40694 ;
  assign n40902 = n40901 ^ n40834 ;
  assign n40903 = n40900 & n40902 ;
  assign n40836 = n40835 ^ n40834 ;
  assign n40695 = n40694 ^ n40691 ;
  assign n40696 = n40694 ^ n38183 ;
  assign n40697 = n40695 & n40696 ;
  assign n40698 = n40697 ^ n38183 ;
  assign n40418 = n40417 ^ n40415 ;
  assign n40142 = n40141 ^ n38374 ;
  assign n40274 = n40273 ^ n40141 ;
  assign n40275 = ~n40142 & ~n40274 ;
  assign n40276 = n40275 ^ n38374 ;
  assign n40310 = n40276 ^ n38466 ;
  assign n40093 = n39739 ^ n39738 ;
  assign n40089 = n39446 ^ n39444 ;
  assign n40088 = n40087 ^ n39446 ;
  assign n40090 = n40089 ^ n40088 ;
  assign n40091 = ~n40086 & n40090 ;
  assign n40092 = n40091 ^ n40089 ;
  assign n40135 = n40093 ^ n40092 ;
  assign n40136 = n38778 & ~n40135 ;
  assign n40137 = n40136 ^ n39446 ;
  assign n40311 = n40310 ^ n40137 ;
  assign n40419 = n40311 ^ x85 ;
  assign n40420 = n40419 ^ n40311 ;
  assign n40421 = n40420 ^ n40415 ;
  assign n40422 = n40418 & n40421 ;
  assign n40423 = n40422 ^ n40419 ;
  assign n40537 = n40423 ^ x84 ;
  assign n40536 = n40533 & n40535 ;
  assign n40568 = n40537 ^ n40536 ;
  assign n40683 = n40568 ^ n40209 ;
  assign n40573 = n40572 ^ n40570 ;
  assign n40574 = n40571 & n40573 ;
  assign n40575 = n40574 ^ n40202 ;
  assign n40684 = n40683 ^ n40575 ;
  assign n40685 = ~n39311 & ~n40684 ;
  assign n40686 = n40685 ^ n40209 ;
  assign n40687 = n40686 ^ n38826 ;
  assign n40831 = n40698 ^ n40687 ;
  assign n40837 = n40831 ^ x294 ;
  assign n40838 = n40837 ^ n40831 ;
  assign n40839 = n40838 ^ n40834 ;
  assign n40840 = ~n40836 & n40839 ;
  assign n40841 = n40840 ^ n40837 ;
  assign n40904 = n40841 ^ x293 ;
  assign n40905 = n40903 & n40904 ;
  assign n40576 = n40575 ^ n40568 ;
  assign n40577 = n40575 ^ n40209 ;
  assign n40578 = ~n40576 & n40577 ;
  assign n40579 = n40578 ^ n40209 ;
  assign n40703 = n40579 ^ n40215 ;
  assign n40312 = n40311 ^ x84 ;
  assign n40424 = ~n40312 & n40423 ;
  assign n40425 = n40424 ^ x84 ;
  assign n40539 = n40425 ^ x83 ;
  assign n40094 = n39741 ^ n39740 ;
  assign n40096 = n40094 ^ n39446 ;
  assign n40095 = n40094 ^ n40093 ;
  assign n40097 = n40096 ^ n40095 ;
  assign n40098 = n40092 & ~n40097 ;
  assign n40099 = n40098 ^ n40096 ;
  assign n40280 = n40099 ^ n39448 ;
  assign n40281 = ~n38773 & n40280 ;
  assign n40282 = n40281 ^ n39448 ;
  assign n40426 = n40282 ^ n38463 ;
  assign n40138 = n40137 ^ n38466 ;
  assign n40277 = n40276 ^ n40137 ;
  assign n40278 = n40138 & n40277 ;
  assign n40279 = n40278 ^ n38466 ;
  assign n40427 = n40426 ^ n40279 ;
  assign n40540 = n40539 ^ n40427 ;
  assign n40538 = ~n40536 & ~n40537 ;
  assign n40566 = n40540 ^ n40538 ;
  assign n40704 = n40703 ^ n40566 ;
  assign n40705 = ~n39313 & n40704 ;
  assign n40706 = n40705 ^ n40215 ;
  assign n40699 = n40698 ^ n40686 ;
  assign n40700 = ~n40687 & ~n40699 ;
  assign n40701 = n40700 ^ n38826 ;
  assign n40702 = n40701 ^ n38836 ;
  assign n40845 = n40706 ^ n40702 ;
  assign n40832 = n40831 ^ x293 ;
  assign n40842 = n40832 & ~n40841 ;
  assign n40843 = n40842 ^ x293 ;
  assign n40844 = n40843 ^ x292 ;
  assign n40906 = n40845 ^ n40844 ;
  assign n40907 = n40905 & ~n40906 ;
  assign n40707 = n40706 ^ n40701 ;
  assign n40708 = ~n40702 & ~n40707 ;
  assign n40709 = n40708 ^ n38836 ;
  assign n40850 = n40709 ^ n38821 ;
  assign n40567 = n40566 ^ n40215 ;
  assign n40580 = n40579 ^ n40566 ;
  assign n40581 = ~n40567 & ~n40580 ;
  assign n40582 = n40581 ^ n40215 ;
  assign n40428 = n40427 ^ n40425 ;
  assign n40283 = n40282 ^ n40279 ;
  assign n40101 = n39450 ^ n39448 ;
  assign n40100 = n40094 ^ n39450 ;
  assign n40102 = n40101 ^ n40100 ;
  assign n40103 = ~n40099 & n40102 ;
  assign n40104 = n40103 ^ n40101 ;
  assign n39757 = n39743 ^ n39742 ;
  assign n40131 = n40104 ^ n39757 ;
  assign n40132 = ~n38922 & ~n40131 ;
  assign n40133 = n40132 ^ n39450 ;
  assign n40284 = n40133 ^ n38463 ;
  assign n40285 = n40284 ^ n40133 ;
  assign n40286 = n40285 ^ n40279 ;
  assign n40287 = ~n40283 & ~n40286 ;
  assign n40288 = n40287 ^ n40284 ;
  assign n40308 = n40288 ^ n38481 ;
  assign n40429 = n40308 ^ x83 ;
  assign n40430 = n40429 ^ n40308 ;
  assign n40431 = n40430 ^ n40425 ;
  assign n40432 = n40428 & n40431 ;
  assign n40433 = n40432 ^ n40429 ;
  assign n40542 = n40433 ^ x82 ;
  assign n40541 = ~n40538 & n40540 ;
  assign n40564 = n40542 ^ n40541 ;
  assign n40565 = n40564 ^ n40191 ;
  assign n40710 = n40582 ^ n40565 ;
  assign n40711 = ~n39315 & ~n40710 ;
  assign n40712 = n40711 ^ n40191 ;
  assign n40851 = n40850 ^ n40712 ;
  assign n40846 = n40845 ^ n40843 ;
  assign n40847 = n40844 & n40846 ;
  assign n40848 = n40847 ^ x292 ;
  assign n40849 = n40848 ^ x291 ;
  assign n40908 = n40851 ^ n40849 ;
  assign n40909 = ~n40907 & n40908 ;
  assign n40852 = n40851 ^ n40848 ;
  assign n40853 = n40849 & n40852 ;
  assign n40854 = n40853 ^ x291 ;
  assign n40910 = n40854 ^ x290 ;
  assign n40713 = n40712 ^ n40709 ;
  assign n40134 = n40133 ^ n38481 ;
  assign n40289 = ~n40134 & ~n40288 ;
  assign n40290 = n40289 ^ n38481 ;
  assign n40436 = n40290 ^ n38459 ;
  assign n39758 = n39757 ^ n39450 ;
  assign n40105 = ~n39758 & ~n40104 ;
  assign n40106 = n40105 ^ n39450 ;
  assign n39755 = n39745 ^ n39744 ;
  assign n39756 = n39755 ^ n39453 ;
  assign n40127 = n40106 ^ n39756 ;
  assign n40128 = ~n38768 & n40127 ;
  assign n40129 = n40128 ^ n39453 ;
  assign n40437 = n40436 ^ n40129 ;
  assign n40544 = n40437 ^ x81 ;
  assign n40309 = n40308 ^ x82 ;
  assign n40434 = n40309 & ~n40433 ;
  assign n40435 = n40434 ^ x82 ;
  assign n40545 = n40544 ^ n40435 ;
  assign n40543 = ~n40541 & n40542 ;
  assign n40586 = n40545 ^ n40543 ;
  assign n40583 = n40582 ^ n40564 ;
  assign n40584 = ~n40565 & ~n40583 ;
  assign n40585 = n40584 ^ n40191 ;
  assign n40587 = n40586 ^ n40585 ;
  assign n40714 = n40587 ^ n40227 ;
  assign n40715 = ~n39318 & ~n40714 ;
  assign n40716 = n40715 ^ n40227 ;
  assign n40717 = n40716 ^ n38821 ;
  assign n40718 = n40717 ^ n40709 ;
  assign n40719 = n40718 ^ n40716 ;
  assign n40720 = ~n40713 & n40719 ;
  assign n40721 = n40720 ^ n40717 ;
  assign n40829 = n40721 ^ n38817 ;
  assign n40911 = n40910 ^ n40829 ;
  assign n40912 = ~n40909 & n40911 ;
  assign n40830 = n40829 ^ x290 ;
  assign n40855 = n40854 ^ n40829 ;
  assign n40856 = n40830 & ~n40855 ;
  assign n40857 = n40856 ^ x290 ;
  assign n40438 = n40437 ^ n40435 ;
  assign n40130 = n40129 ^ n38459 ;
  assign n40291 = n40290 ^ n40129 ;
  assign n40292 = ~n40130 & n40291 ;
  assign n40293 = n40292 ^ n38459 ;
  assign n40107 = n40106 ^ n39755 ;
  assign n40108 = ~n39756 & n40107 ;
  assign n40109 = n40108 ^ n39453 ;
  assign n39753 = n39746 ^ n39721 ;
  assign n39754 = n39753 ^ n39437 ;
  assign n40123 = n40109 ^ n39754 ;
  assign n40124 = ~n38933 & n40123 ;
  assign n40125 = n40124 ^ n39437 ;
  assign n40126 = n40125 ^ n38492 ;
  assign n40306 = n40293 ^ n40126 ;
  assign n40439 = n40306 ^ x81 ;
  assign n40440 = n40439 ^ n40306 ;
  assign n40441 = n40440 ^ n40435 ;
  assign n40442 = n40438 & n40441 ;
  assign n40443 = n40442 ^ n40439 ;
  assign n40547 = n40443 ^ x80 ;
  assign n40546 = ~n40543 & n40545 ;
  assign n40562 = n40547 ^ n40546 ;
  assign n40589 = n40562 ^ n40227 ;
  assign n40588 = n40585 ^ n40562 ;
  assign n40590 = n40589 ^ n40588 ;
  assign n40591 = ~n40587 & n40590 ;
  assign n40592 = n40591 ^ n40589 ;
  assign n40679 = n40592 ^ n40187 ;
  assign n40680 = n39320 & n40679 ;
  assign n40681 = n40680 ^ n40187 ;
  assign n40723 = n40681 ^ n38817 ;
  assign n40722 = n40716 ^ n40681 ;
  assign n40724 = n40723 ^ n40722 ;
  assign n40725 = ~n40721 & ~n40724 ;
  assign n40726 = n40725 ^ n40723 ;
  assign n40827 = n40726 ^ n38389 ;
  assign n40828 = n40827 ^ x289 ;
  assign n40913 = n40857 ^ n40828 ;
  assign n40914 = n40912 & ~n40913 ;
  assign n40682 = n40681 ^ n38389 ;
  assign n40727 = ~n40682 & n40726 ;
  assign n40728 = n40727 ^ n38389 ;
  assign n40563 = n40562 ^ n40187 ;
  assign n40593 = ~n40563 & n40592 ;
  assign n40594 = n40593 ^ n40187 ;
  assign n40307 = n40306 ^ x80 ;
  assign n40444 = ~n40307 & n40443 ;
  assign n40445 = n40444 ^ x80 ;
  assign n40549 = n40445 ^ x95 ;
  assign n40294 = n40293 ^ n40125 ;
  assign n40295 = ~n40126 & ~n40294 ;
  assign n40296 = n40295 ^ n38492 ;
  assign n40303 = n40296 ^ n38423 ;
  assign n40110 = n40109 ^ n39753 ;
  assign n40111 = ~n39754 & ~n40110 ;
  assign n40112 = n40111 ^ n39437 ;
  assign n39751 = n39747 ^ n39720 ;
  assign n39752 = n39751 ^ n39469 ;
  assign n40119 = n40112 ^ n39752 ;
  assign n40120 = n38939 & ~n40119 ;
  assign n40121 = n40120 ^ n39469 ;
  assign n40304 = n40303 ^ n40121 ;
  assign n40550 = n40549 ^ n40304 ;
  assign n40548 = n40546 & n40547 ;
  assign n40560 = n40550 ^ n40548 ;
  assign n40561 = n40560 ^ n40183 ;
  assign n40675 = n40594 ^ n40561 ;
  assign n40676 = n39307 & ~n40675 ;
  assign n40677 = n40676 ^ n40183 ;
  assign n40678 = n40677 ^ n38386 ;
  assign n40861 = n40728 ^ n40678 ;
  assign n40915 = n40861 ^ x288 ;
  assign n40858 = n40857 ^ n40827 ;
  assign n40859 = ~n40828 & n40858 ;
  assign n40860 = n40859 ^ x289 ;
  assign n40916 = n40915 ^ n40860 ;
  assign n40917 = ~n40914 & n40916 ;
  assign n40862 = n40861 ^ n40860 ;
  assign n40729 = n40728 ^ n40677 ;
  assign n40730 = ~n40678 & ~n40729 ;
  assign n40731 = n40730 ^ n38386 ;
  assign n40595 = n40594 ^ n40560 ;
  assign n40596 = n40561 & n40595 ;
  assign n40597 = n40596 ^ n40183 ;
  assign n40670 = n40597 ^ n40178 ;
  assign n40305 = n40304 ^ x95 ;
  assign n40446 = n40445 ^ n40304 ;
  assign n40447 = n40305 & ~n40446 ;
  assign n40448 = n40447 ^ x95 ;
  assign n40122 = n40121 ^ n38423 ;
  assign n40297 = n40296 ^ n40121 ;
  assign n40298 = ~n40122 & n40297 ;
  assign n40299 = n40298 ^ n38423 ;
  assign n40300 = n40299 ^ n38504 ;
  assign n40113 = n40112 ^ n39751 ;
  assign n40114 = ~n39752 & n40113 ;
  assign n40115 = n40114 ^ n39469 ;
  assign n39749 = n39748 ^ n39719 ;
  assign n39750 = n39749 ^ n39478 ;
  assign n40116 = n40115 ^ n39750 ;
  assign n40117 = n38764 & n40116 ;
  assign n40118 = n40117 ^ n39478 ;
  assign n40301 = n40300 ^ n40118 ;
  assign n40302 = n40301 ^ x94 ;
  assign n40552 = n40448 ^ n40302 ;
  assign n40551 = ~n40548 & n40550 ;
  assign n40558 = n40552 ^ n40551 ;
  assign n40671 = n40670 ^ n40558 ;
  assign n40672 = ~n39374 & n40671 ;
  assign n40673 = n40672 ^ n40178 ;
  assign n40674 = n40673 ^ n38862 ;
  assign n40825 = n40731 ^ n40674 ;
  assign n40863 = n40825 ^ x288 ;
  assign n40864 = n40863 ^ n40825 ;
  assign n40865 = n40864 ^ n40860 ;
  assign n40866 = n40862 & n40865 ;
  assign n40867 = n40866 ^ n40863 ;
  assign n40918 = n40867 ^ x303 ;
  assign n40919 = n40917 & n40918 ;
  assign n40732 = n40731 ^ n40673 ;
  assign n40733 = n40674 & n40732 ;
  assign n40734 = n40733 ^ n38862 ;
  assign n40559 = n40558 ^ n40178 ;
  assign n40598 = n40597 ^ n40558 ;
  assign n40599 = n40559 & ~n40598 ;
  assign n40600 = n40599 ^ n40178 ;
  assign n40553 = ~n40551 & ~n40552 ;
  assign n40462 = n39970 ^ n39968 ;
  assign n40456 = n40115 ^ n39749 ;
  assign n40457 = n39486 ^ n39478 ;
  assign n40458 = n40457 ^ n39486 ;
  assign n40459 = n40458 ^ n39749 ;
  assign n40460 = ~n40456 & n40459 ;
  assign n40461 = n40460 ^ n40457 ;
  assign n40463 = n40462 ^ n40461 ;
  assign n40464 = n38956 & ~n40463 ;
  assign n40465 = n40464 ^ n39486 ;
  assign n40452 = n40299 ^ n40118 ;
  assign n40453 = n40300 & n40452 ;
  assign n40454 = n40453 ^ n38504 ;
  assign n40455 = n40454 ^ n38508 ;
  assign n40466 = n40465 ^ n40455 ;
  assign n40489 = n40466 ^ x93 ;
  assign n40449 = n40448 ^ n40301 ;
  assign n40450 = n40302 & ~n40449 ;
  assign n40451 = n40450 ^ x94 ;
  assign n40490 = n40489 ^ n40451 ;
  assign n40556 = n40553 ^ n40490 ;
  assign n40557 = n40556 ^ n40174 ;
  assign n40666 = n40600 ^ n40557 ;
  assign n40667 = ~n39376 & n40666 ;
  assign n40668 = n40667 ^ n40174 ;
  assign n40669 = n40668 ^ n38866 ;
  assign n40870 = n40734 ^ n40669 ;
  assign n40920 = n40870 ^ x302 ;
  assign n40826 = n40825 ^ x303 ;
  assign n40868 = ~n40826 & n40867 ;
  assign n40869 = n40868 ^ x303 ;
  assign n40921 = n40920 ^ n40869 ;
  assign n40922 = n40919 & ~n40921 ;
  assign n40871 = n40870 ^ n40869 ;
  assign n40735 = n40734 ^ n40668 ;
  assign n40736 = n40669 & n40735 ;
  assign n40737 = n40736 ^ n38866 ;
  assign n40554 = ~n40490 & ~n40553 ;
  assign n40467 = n40466 ^ n40451 ;
  assign n40473 = n39972 ^ n39971 ;
  assign n40475 = n40473 ^ n39486 ;
  assign n40474 = n40473 ^ n40462 ;
  assign n40476 = n40475 ^ n40474 ;
  assign n40477 = n40461 & ~n40476 ;
  assign n40478 = n40477 ^ n40475 ;
  assign n40479 = n40478 ^ n39494 ;
  assign n40480 = n38969 & n40479 ;
  assign n40481 = n40480 ^ n39494 ;
  assign n40468 = n40465 ^ n40454 ;
  assign n40469 = n40465 ^ n38508 ;
  assign n40470 = n40468 & n40469 ;
  assign n40471 = n40470 ^ n38508 ;
  assign n40472 = n40471 ^ n38452 ;
  assign n40482 = n40481 ^ n40472 ;
  assign n40483 = n40482 ^ x93 ;
  assign n40484 = n40483 ^ n40451 ;
  assign n40485 = n40484 ^ n40482 ;
  assign n40486 = n40467 & n40485 ;
  assign n40487 = n40486 ^ n40483 ;
  assign n40488 = n40487 ^ x92 ;
  assign n40555 = n40554 ^ n40488 ;
  assign n40661 = n40555 ^ n40245 ;
  assign n40601 = n40600 ^ n40556 ;
  assign n40602 = n40557 & n40601 ;
  assign n40603 = n40602 ^ n40174 ;
  assign n40662 = n40661 ^ n40603 ;
  assign n40663 = ~n39378 & ~n40662 ;
  assign n40664 = n40663 ^ n40245 ;
  assign n40665 = n40664 ^ n38810 ;
  assign n40823 = n40737 ^ n40665 ;
  assign n40872 = n40823 ^ x302 ;
  assign n40873 = n40872 ^ n40823 ;
  assign n40874 = n40873 ^ n40869 ;
  assign n40875 = ~n40871 & n40874 ;
  assign n40876 = n40875 ^ n40872 ;
  assign n40923 = n40876 ^ x301 ;
  assign n40924 = ~n40922 & ~n40923 ;
  assign n40604 = n40603 ^ n40555 ;
  assign n40605 = n40603 ^ n40245 ;
  assign n40606 = n40604 & ~n40605 ;
  assign n40607 = n40606 ^ n40245 ;
  assign n40742 = n40607 ^ n40169 ;
  assign n40627 = ~n40488 & ~n40554 ;
  assign n40619 = n40473 ^ n39494 ;
  assign n40620 = n40478 & n40619 ;
  assign n40621 = n40620 ^ n39494 ;
  assign n40617 = n39974 ^ n39973 ;
  assign n40618 = n40617 ^ n39502 ;
  assign n40622 = n40621 ^ n40618 ;
  assign n40623 = ~n38982 & ~n40622 ;
  assign n40624 = n40623 ^ n39502 ;
  assign n40612 = n40481 ^ n40471 ;
  assign n40613 = n40481 ^ n38452 ;
  assign n40614 = n40612 & n40613 ;
  assign n40615 = n40614 ^ n38452 ;
  assign n40616 = n40615 ^ n38448 ;
  assign n40625 = n40624 ^ n40616 ;
  assign n40608 = n40482 ^ x92 ;
  assign n40609 = ~n40487 & n40608 ;
  assign n40610 = n40609 ^ x92 ;
  assign n40611 = n40610 ^ x91 ;
  assign n40626 = n40625 ^ n40611 ;
  assign n40628 = n40627 ^ n40626 ;
  assign n40743 = n40742 ^ n40628 ;
  assign n40744 = n39380 & ~n40743 ;
  assign n40745 = n40744 ^ n40169 ;
  assign n40738 = n40737 ^ n40664 ;
  assign n40739 = n40665 & n40738 ;
  assign n40740 = n40739 ^ n38810 ;
  assign n40741 = n40740 ^ n38805 ;
  assign n40879 = n40745 ^ n40741 ;
  assign n40898 = n40879 ^ x300 ;
  assign n40824 = n40823 ^ x301 ;
  assign n40877 = ~n40824 & n40876 ;
  assign n40878 = n40877 ^ x301 ;
  assign n40899 = n40898 ^ n40878 ;
  assign n40949 = n40924 ^ n40899 ;
  assign n41051 = n40949 ^ n40688 ;
  assign n40950 = n40688 & n40949 ;
  assign n41052 = n40950 ^ n40692 ;
  assign n40925 = n40899 & n40924 ;
  assign n40880 = n40879 ^ n40878 ;
  assign n40629 = n40628 ^ n40607 ;
  assign n40651 = ~n40626 & ~n40627 ;
  assign n40635 = n40624 ^ n40615 ;
  assign n40639 = n39976 ^ n39975 ;
  assign n40636 = n40621 ^ n39502 ;
  assign n40637 = n40618 & n40636 ;
  assign n40638 = n40637 ^ n39502 ;
  assign n40640 = n40639 ^ n40638 ;
  assign n40641 = n40640 ^ n39509 ;
  assign n40642 = ~n38995 & n40641 ;
  assign n40643 = n40642 ^ n39509 ;
  assign n40644 = n40643 ^ n38448 ;
  assign n40645 = n40644 ^ n40643 ;
  assign n40646 = n40645 ^ n40615 ;
  assign n40647 = ~n40635 & n40646 ;
  assign n40648 = n40647 ^ n40644 ;
  assign n40649 = n40648 ^ n38533 ;
  assign n40630 = n40625 ^ n40610 ;
  assign n40631 = n40625 ^ x91 ;
  assign n40632 = n40630 & ~n40631 ;
  assign n40633 = n40632 ^ x91 ;
  assign n40634 = n40633 ^ x90 ;
  assign n40650 = n40649 ^ n40634 ;
  assign n40652 = n40651 ^ n40650 ;
  assign n40653 = n40652 ^ n40169 ;
  assign n40654 = n40653 ^ n40652 ;
  assign n40655 = n40654 ^ n40607 ;
  assign n40656 = n40629 & n40655 ;
  assign n40657 = n40656 ^ n40653 ;
  assign n40658 = n40657 ^ n40165 ;
  assign n40659 = n39382 & ~n40658 ;
  assign n40660 = n40659 ^ n40165 ;
  assign n40820 = n40660 ^ n38884 ;
  assign n40746 = n40745 ^ n40740 ;
  assign n40747 = n40741 & ~n40746 ;
  assign n40748 = n40747 ^ n38805 ;
  assign n40821 = n40820 ^ n40748 ;
  assign n40881 = n40821 ^ x300 ;
  assign n40882 = n40881 ^ n40878 ;
  assign n40883 = n40882 ^ n40821 ;
  assign n40884 = ~n40880 & n40883 ;
  assign n40885 = n40884 ^ n40881 ;
  assign n40897 = n40885 ^ x299 ;
  assign n40951 = n40925 ^ n40897 ;
  assign n41053 = n41052 ^ n40951 ;
  assign n41054 = n41051 & ~n41053 ;
  assign n40952 = n40951 ^ n40950 ;
  assign n40953 = n40951 ^ n40692 ;
  assign n40954 = ~n40952 & ~n40953 ;
  assign n40955 = n40954 ^ n40692 ;
  assign n41055 = n40955 ^ n40684 ;
  assign n40926 = n40897 & ~n40925 ;
  assign n40749 = n40748 ^ n40660 ;
  assign n40750 = n40748 ^ n38884 ;
  assign n40751 = n40749 & n40750 ;
  assign n40752 = n40751 ^ n38884 ;
  assign n40889 = n40752 ^ n38800 ;
  assign n40777 = ~n40650 & ~n40651 ;
  assign n40771 = n40643 ^ n38533 ;
  assign n40772 = ~n40648 & ~n40771 ;
  assign n40773 = n40772 ^ n38533 ;
  assign n40761 = n39979 ^ n39977 ;
  assign n40762 = n40761 ^ n39509 ;
  assign n40763 = n40762 ^ n40638 ;
  assign n40764 = n40763 ^ n40761 ;
  assign n40765 = n40640 & n40764 ;
  assign n40766 = n40765 ^ n40762 ;
  assign n40767 = n40766 ^ n39516 ;
  assign n40768 = n39009 & ~n40767 ;
  assign n40769 = n40768 ^ n39516 ;
  assign n40770 = n40769 ^ n38543 ;
  assign n40774 = n40773 ^ n40770 ;
  assign n40775 = n40774 ^ x89 ;
  assign n40757 = n40649 ^ n40633 ;
  assign n40758 = n40649 ^ x90 ;
  assign n40759 = ~n40757 & n40758 ;
  assign n40760 = n40759 ^ x90 ;
  assign n40776 = n40775 ^ n40760 ;
  assign n40778 = n40777 ^ n40776 ;
  assign n40753 = n40652 ^ n40165 ;
  assign n40754 = ~n40657 & ~n40753 ;
  assign n40755 = n40754 ^ n40165 ;
  assign n40756 = n40755 ^ n40161 ;
  assign n40779 = n40778 ^ n40756 ;
  assign n40780 = ~n39384 & ~n40779 ;
  assign n40781 = n40780 ^ n40161 ;
  assign n40890 = n40889 ^ n40781 ;
  assign n40822 = n40821 ^ x299 ;
  assign n40886 = ~n40822 & n40885 ;
  assign n40887 = n40886 ^ x299 ;
  assign n40888 = n40887 ^ x298 ;
  assign n40896 = n40890 ^ n40888 ;
  assign n40956 = n40926 ^ n40896 ;
  assign n41056 = n41055 ^ n40956 ;
  assign n41057 = n41054 & n41056 ;
  assign n40957 = n40956 ^ n40955 ;
  assign n40927 = n40896 & ~n40926 ;
  assign n40891 = n40890 ^ n40887 ;
  assign n40892 = n40888 & ~n40891 ;
  assign n40893 = n40892 ^ x298 ;
  assign n40894 = n40893 ^ x297 ;
  assign n40782 = n40781 ^ n40752 ;
  assign n40806 = n40778 ^ n40755 ;
  assign n40807 = n40778 ^ n40161 ;
  assign n40808 = ~n40806 & n40807 ;
  assign n40809 = n40808 ^ n40161 ;
  assign n40810 = n40809 ^ n40157 ;
  assign n40800 = n40761 ^ n39516 ;
  assign n40801 = n40766 & n40800 ;
  assign n40797 = n39982 ^ n39980 ;
  assign n40798 = n40797 ^ n39523 ;
  assign n40799 = n40798 ^ n40761 ;
  assign n40802 = n40801 ^ n40799 ;
  assign n40803 = ~n39207 & ~n40802 ;
  assign n40793 = n38636 ^ n38543 ;
  assign n40794 = n40793 ^ n39523 ;
  assign n40795 = n40794 ^ x88 ;
  assign n40790 = n40773 ^ n40769 ;
  assign n40791 = n40773 ^ n38543 ;
  assign n40792 = n40790 & n40791 ;
  assign n40796 = n40795 ^ n40792 ;
  assign n40804 = n40803 ^ n40796 ;
  assign n40783 = n40777 ^ n40774 ;
  assign n40785 = n40774 ^ n40760 ;
  assign n40788 = ~n40783 & n40785 ;
  assign n40786 = n40785 ^ n40777 ;
  assign n40787 = ~x89 & n40786 ;
  assign n40789 = n40788 ^ n40787 ;
  assign n40805 = n40804 ^ n40789 ;
  assign n40811 = n40810 ^ n40805 ;
  assign n40812 = n39386 & n40811 ;
  assign n40813 = n40812 ^ n40157 ;
  assign n40814 = n40813 ^ n38800 ;
  assign n40815 = n40814 ^ n40813 ;
  assign n40816 = n40815 ^ n40752 ;
  assign n40817 = n40782 & ~n40816 ;
  assign n40818 = n40817 ^ n40814 ;
  assign n40819 = n40818 ^ n38795 ;
  assign n40895 = n40894 ^ n40819 ;
  assign n40958 = n40927 ^ n40895 ;
  assign n40959 = n40958 ^ n40684 ;
  assign n40960 = n40959 ^ n40958 ;
  assign n40961 = n40960 ^ n40955 ;
  assign n40962 = ~n40957 & ~n40961 ;
  assign n40963 = n40962 ^ n40959 ;
  assign n41058 = n40963 ^ n40704 ;
  assign n41059 = ~n41057 & n41058 ;
  assign n40940 = n40491 ^ n40153 ;
  assign n40936 = n40809 ^ n40805 ;
  assign n40937 = n40805 ^ n40157 ;
  assign n40938 = n40936 & ~n40937 ;
  assign n40939 = n40938 ^ n40157 ;
  assign n40941 = n40940 ^ n40939 ;
  assign n40942 = n39372 & n40941 ;
  assign n40943 = n40942 ^ n40153 ;
  assign n40932 = n40813 ^ n38795 ;
  assign n40933 = ~n40818 & n40932 ;
  assign n40934 = n40933 ^ n38795 ;
  assign n40935 = n40934 ^ n38791 ;
  assign n40944 = n40943 ^ n40935 ;
  assign n40945 = n40944 ^ x296 ;
  assign n40929 = n40893 ^ n40819 ;
  assign n40930 = n40894 & n40929 ;
  assign n40931 = n40930 ^ x297 ;
  assign n40946 = n40945 ^ n40931 ;
  assign n40928 = n40895 & ~n40927 ;
  assign n40947 = n40946 ^ n40928 ;
  assign n40965 = n40947 ^ n40704 ;
  assign n40964 = n40958 ^ n40947 ;
  assign n40966 = n40965 ^ n40964 ;
  assign n40967 = ~n40963 & ~n40966 ;
  assign n40968 = n40967 ^ n40965 ;
  assign n41060 = n40968 ^ n40710 ;
  assign n41061 = ~n41059 & ~n41060 ;
  assign n40994 = n40928 & ~n40946 ;
  assign n40972 = n40944 ^ n40931 ;
  assign n40973 = n40943 ^ n40934 ;
  assign n40976 = n40939 ^ n40491 ;
  assign n40977 = ~n40940 & ~n40976 ;
  assign n40978 = n40977 ^ n40153 ;
  assign n40974 = n40493 ^ n40491 ;
  assign n40975 = n40974 ^ n40148 ;
  assign n40979 = n40978 ^ n40975 ;
  assign n40980 = n39440 & n40979 ;
  assign n40981 = n40980 ^ n40148 ;
  assign n40982 = n40981 ^ n38791 ;
  assign n40983 = n40982 ^ n40934 ;
  assign n40984 = n40983 ^ n40981 ;
  assign n40985 = n40973 & n40984 ;
  assign n40986 = n40985 ^ n40982 ;
  assign n40987 = n40986 ^ n38901 ;
  assign n40988 = n40987 ^ x296 ;
  assign n40989 = n40988 ^ n40931 ;
  assign n40990 = n40989 ^ n40987 ;
  assign n40991 = ~n40972 & n40990 ;
  assign n40992 = n40991 ^ n40988 ;
  assign n40993 = n40992 ^ x311 ;
  assign n40995 = n40994 ^ n40993 ;
  assign n40948 = n40947 ^ n40710 ;
  assign n40969 = n40948 & n40968 ;
  assign n40970 = n40969 ^ n40710 ;
  assign n40971 = n40970 ^ n40714 ;
  assign n41062 = n40995 ^ n40971 ;
  assign n41063 = n41061 & ~n41062 ;
  assign n41021 = n40993 & ~n40994 ;
  assign n40999 = n40978 ^ n40974 ;
  assign n41000 = n40496 ^ n40494 ;
  assign n41001 = n41000 ^ n40148 ;
  assign n41002 = n41001 ^ n40974 ;
  assign n41003 = n41002 ^ n41000 ;
  assign n41004 = ~n40999 & n41003 ;
  assign n41005 = n41004 ^ n41001 ;
  assign n41006 = n41005 ^ n40144 ;
  assign n41007 = n39442 & ~n41006 ;
  assign n41008 = n41007 ^ n40144 ;
  assign n41010 = n41008 ^ n38901 ;
  assign n41009 = n41008 ^ n40981 ;
  assign n41011 = n41010 ^ n41009 ;
  assign n41012 = n40986 & ~n41011 ;
  assign n41013 = n41012 ^ n41010 ;
  assign n41014 = n41013 ^ n38786 ;
  assign n41016 = n41014 ^ x311 ;
  assign n41015 = n41014 ^ n40987 ;
  assign n41017 = n41016 ^ n41015 ;
  assign n41018 = ~n40992 & n41017 ;
  assign n41019 = n41018 ^ n41016 ;
  assign n41020 = n41019 ^ x310 ;
  assign n41022 = n41021 ^ n41020 ;
  assign n41064 = n41022 ^ n40679 ;
  assign n40996 = n40995 ^ n40970 ;
  assign n40997 = n40971 & n40996 ;
  assign n40998 = n40997 ^ n40714 ;
  assign n41065 = n41064 ^ n40998 ;
  assign n41066 = n41063 & ~n41065 ;
  assign n41023 = n41022 ^ n40998 ;
  assign n41043 = n41020 & ~n41021 ;
  assign n41030 = n41000 ^ n40144 ;
  assign n41031 = n41005 & ~n41030 ;
  assign n41029 = n40144 ^ n40139 ;
  assign n41032 = n41031 ^ n41029 ;
  assign n41028 = n40498 ^ n40497 ;
  assign n41033 = n41032 ^ n41028 ;
  assign n41034 = ~n39444 & ~n41033 ;
  assign n41035 = n41034 ^ n40139 ;
  assign n41024 = n41008 ^ n38786 ;
  assign n41025 = n41013 & n41024 ;
  assign n41026 = n41025 ^ n38786 ;
  assign n41027 = n41026 ^ n38782 ;
  assign n41036 = n41035 ^ n41027 ;
  assign n41038 = n41036 ^ x310 ;
  assign n41037 = n41036 ^ n41014 ;
  assign n41039 = n41038 ^ n41037 ;
  assign n41040 = n41019 & ~n41039 ;
  assign n41041 = n41040 ^ n41038 ;
  assign n41042 = n41041 ^ x309 ;
  assign n41044 = n41043 ^ n41042 ;
  assign n41045 = n41044 ^ n40679 ;
  assign n41046 = n41045 ^ n40998 ;
  assign n41047 = n41046 ^ n41044 ;
  assign n41048 = ~n41023 & ~n41047 ;
  assign n41049 = n41048 ^ n41045 ;
  assign n41050 = n41049 ^ n40675 ;
  assign n41067 = n41066 ^ n41050 ;
  assign n41068 = n41065 ^ n41063 ;
  assign n41069 = n41062 ^ n41061 ;
  assign n41070 = n41060 ^ n41059 ;
  assign n41071 = n41058 ^ n41057 ;
  assign n41072 = n41056 ^ n41054 ;
  assign n41073 = n41053 ^ n41051 ;
  assign n41285 = ~n41050 & ~n41066 ;
  assign n41174 = n41042 & n41043 ;
  assign n41092 = n41035 ^ n41026 ;
  assign n41093 = n41035 ^ n38782 ;
  assign n41094 = n41092 & ~n41093 ;
  assign n41095 = n41094 ^ n38782 ;
  assign n41074 = n40500 ^ n40499 ;
  assign n41087 = n41074 ^ n40135 ;
  assign n41075 = n41028 ^ n40139 ;
  assign n41076 = ~n41032 & ~n41075 ;
  assign n41077 = n41076 ^ n40139 ;
  assign n41088 = n41087 ^ n41077 ;
  assign n41089 = ~n39446 & ~n41088 ;
  assign n41090 = n41089 ^ n40135 ;
  assign n41091 = n41090 ^ n38778 ;
  assign n41128 = n41095 ^ n41091 ;
  assign n41131 = n41128 ^ x309 ;
  assign n41130 = n41128 ^ n41036 ;
  assign n41132 = n41131 ^ n41130 ;
  assign n41133 = n41041 & ~n41132 ;
  assign n41134 = n41133 ^ n41131 ;
  assign n41173 = n41134 ^ x308 ;
  assign n41211 = n41174 ^ n41173 ;
  assign n41286 = n41211 ^ n40671 ;
  assign n41208 = n41044 ^ n40675 ;
  assign n41209 = ~n41049 & ~n41208 ;
  assign n41210 = n41209 ^ n40675 ;
  assign n41287 = n41286 ^ n41210 ;
  assign n41288 = n41285 & n41287 ;
  assign n41212 = n41211 ^ n41210 ;
  assign n41175 = ~n41173 & ~n41174 ;
  assign n41082 = n40503 ^ n40501 ;
  assign n41083 = n41082 ^ n40280 ;
  assign n41078 = n41077 ^ n41074 ;
  assign n41079 = n41077 ^ n40135 ;
  assign n41080 = ~n41078 & n41079 ;
  assign n41081 = n41080 ^ n40135 ;
  assign n41084 = n41083 ^ n41081 ;
  assign n41085 = ~n39448 & n41084 ;
  assign n41086 = n41085 ^ n40280 ;
  assign n41137 = n41086 ^ n38773 ;
  assign n41096 = n41095 ^ n41090 ;
  assign n41097 = ~n41091 & n41096 ;
  assign n41098 = n41097 ^ n38778 ;
  assign n41138 = n41137 ^ n41098 ;
  assign n41171 = n41138 ^ x307 ;
  assign n41129 = n41128 ^ x308 ;
  assign n41135 = ~n41129 & n41134 ;
  assign n41136 = n41135 ^ x308 ;
  assign n41172 = n41171 ^ n41136 ;
  assign n41206 = n41175 ^ n41172 ;
  assign n41213 = n41206 ^ n40671 ;
  assign n41214 = n41213 ^ n41210 ;
  assign n41215 = n41214 ^ n41206 ;
  assign n41216 = ~n41212 & ~n41215 ;
  assign n41217 = n41216 ^ n41213 ;
  assign n41289 = n41217 ^ n40666 ;
  assign n41290 = n41288 & n41289 ;
  assign n41207 = n41206 ^ n40666 ;
  assign n41218 = n41207 & ~n41217 ;
  assign n41219 = n41218 ^ n40666 ;
  assign n41291 = n41219 ^ n40662 ;
  assign n41176 = ~n41172 & n41175 ;
  assign n41139 = n41138 ^ n41136 ;
  assign n41099 = n41098 ^ n41086 ;
  assign n41100 = n41098 ^ n38773 ;
  assign n41101 = ~n41099 & ~n41100 ;
  assign n41102 = n41101 ^ n38773 ;
  assign n41125 = n41102 ^ n38922 ;
  assign n41105 = n41082 ^ n41081 ;
  assign n41106 = ~n41083 & ~n41105 ;
  assign n41104 = n40280 ^ n40131 ;
  assign n41107 = n41106 ^ n41104 ;
  assign n41103 = n40506 ^ n40504 ;
  assign n41108 = n41107 ^ n41103 ;
  assign n41109 = n39450 & n41108 ;
  assign n41110 = n41109 ^ n40131 ;
  assign n41126 = n41125 ^ n41110 ;
  assign n41140 = n41126 ^ x307 ;
  assign n41141 = n41140 ^ n41136 ;
  assign n41142 = n41141 ^ n41126 ;
  assign n41143 = n41139 & n41142 ;
  assign n41144 = n41143 ^ n41140 ;
  assign n41170 = n41144 ^ x306 ;
  assign n41205 = n41176 ^ n41170 ;
  assign n41292 = n41291 ^ n41205 ;
  assign n41293 = ~n41290 & n41292 ;
  assign n41220 = n41219 ^ n41205 ;
  assign n41177 = ~n41170 & n41176 ;
  assign n41127 = n41126 ^ x306 ;
  assign n41145 = ~n41127 & n41144 ;
  assign n41146 = n41145 ^ x306 ;
  assign n41168 = n41146 ^ x305 ;
  assign n41118 = n41103 ^ n40131 ;
  assign n41119 = ~n41107 & n41118 ;
  assign n41120 = n41119 ^ n40131 ;
  assign n41116 = n40509 ^ n40507 ;
  assign n41117 = n41116 ^ n40127 ;
  assign n41121 = n41120 ^ n41117 ;
  assign n41122 = n39453 & ~n41121 ;
  assign n41123 = n41122 ^ n40127 ;
  assign n41111 = n41110 ^ n41102 ;
  assign n41112 = n41110 ^ n38922 ;
  assign n41113 = ~n41111 & n41112 ;
  assign n41114 = n41113 ^ n38922 ;
  assign n41115 = n41114 ^ n38768 ;
  assign n41124 = n41123 ^ n41115 ;
  assign n41169 = n41168 ^ n41124 ;
  assign n41203 = n41177 ^ n41169 ;
  assign n41221 = n41203 ^ n40662 ;
  assign n41222 = n41221 ^ n41205 ;
  assign n41223 = n41222 ^ n41203 ;
  assign n41224 = ~n41220 & ~n41223 ;
  assign n41225 = n41224 ^ n41221 ;
  assign n41294 = n41225 ^ n40743 ;
  assign n41295 = ~n41293 & ~n41294 ;
  assign n41204 = n41203 ^ n40743 ;
  assign n41226 = n41204 & ~n41225 ;
  assign n41227 = n41226 ^ n40743 ;
  assign n41296 = n41227 ^ n40658 ;
  assign n41178 = n41169 & n41177 ;
  assign n41147 = n41146 ^ n41124 ;
  assign n41157 = n40511 ^ n40510 ;
  assign n41154 = n41120 ^ n40127 ;
  assign n41155 = n41117 & ~n41154 ;
  assign n41153 = n40127 ^ n40123 ;
  assign n41156 = n41155 ^ n41153 ;
  assign n41158 = n41157 ^ n41156 ;
  assign n41159 = ~n39437 & ~n41158 ;
  assign n41160 = n41159 ^ n40123 ;
  assign n41148 = n41123 ^ n41114 ;
  assign n41149 = n41123 ^ n38768 ;
  assign n41150 = n41148 & ~n41149 ;
  assign n41151 = n41150 ^ n38768 ;
  assign n41152 = n41151 ^ n38933 ;
  assign n41161 = n41160 ^ n41152 ;
  assign n41162 = n41161 ^ x305 ;
  assign n41163 = n41162 ^ n41124 ;
  assign n41164 = n41163 ^ n41161 ;
  assign n41165 = ~n41147 & n41164 ;
  assign n41166 = n41165 ^ n41162 ;
  assign n41167 = n41166 ^ x304 ;
  assign n41202 = n41178 ^ n41167 ;
  assign n41297 = n41296 ^ n41202 ;
  assign n41298 = ~n41295 & ~n41297 ;
  assign n41228 = n41227 ^ n41202 ;
  assign n41186 = n41157 ^ n40123 ;
  assign n41187 = n41156 & ~n41186 ;
  assign n41188 = n41187 ^ n40123 ;
  assign n41184 = n40514 ^ n40512 ;
  assign n41185 = n41184 ^ n40119 ;
  assign n41189 = n41188 ^ n41185 ;
  assign n41190 = ~n39469 & ~n41189 ;
  assign n41191 = n41190 ^ n40119 ;
  assign n41192 = n41191 ^ n38939 ;
  assign n41180 = n41160 ^ n41151 ;
  assign n41181 = n41160 ^ n38933 ;
  assign n41182 = n41180 & ~n41181 ;
  assign n41183 = n41182 ^ n38933 ;
  assign n41193 = n41192 ^ n41183 ;
  assign n41195 = n41193 ^ x304 ;
  assign n41194 = n41193 ^ n41161 ;
  assign n41196 = n41195 ^ n41194 ;
  assign n41197 = ~n41166 & n41196 ;
  assign n41198 = n41197 ^ n41195 ;
  assign n41199 = n41198 ^ x319 ;
  assign n41179 = ~n41167 & ~n41178 ;
  assign n41200 = n41199 ^ n41179 ;
  assign n41229 = n41200 ^ n40658 ;
  assign n41230 = n41229 ^ n41202 ;
  assign n41231 = n41230 ^ n41200 ;
  assign n41232 = n41228 & ~n41231 ;
  assign n41233 = n41232 ^ n41229 ;
  assign n41299 = n41233 ^ n40779 ;
  assign n41300 = ~n41298 & ~n41299 ;
  assign n41256 = n41179 & ~n41199 ;
  assign n41244 = n40517 ^ n40515 ;
  assign n41241 = n41188 ^ n40119 ;
  assign n41242 = ~n41185 & ~n41241 ;
  assign n41243 = n41242 ^ n40119 ;
  assign n41245 = n41244 ^ n41243 ;
  assign n41246 = n41245 ^ n40116 ;
  assign n41247 = ~n39478 & n41246 ;
  assign n41248 = n41247 ^ n40116 ;
  assign n41237 = n41191 ^ n41183 ;
  assign n41238 = ~n41192 & ~n41237 ;
  assign n41239 = n41238 ^ n38939 ;
  assign n41240 = n41239 ^ n38764 ;
  assign n41249 = n41248 ^ n41240 ;
  assign n41251 = n41249 ^ x319 ;
  assign n41250 = n41249 ^ n41193 ;
  assign n41252 = n41251 ^ n41250 ;
  assign n41253 = ~n41198 & n41252 ;
  assign n41254 = n41253 ^ n41251 ;
  assign n41255 = n41254 ^ x318 ;
  assign n41257 = n41256 ^ n41255 ;
  assign n41201 = n41200 ^ n40779 ;
  assign n41234 = n41201 & ~n41233 ;
  assign n41235 = n41234 ^ n40779 ;
  assign n41236 = n41235 ^ n40811 ;
  assign n41301 = n41257 ^ n41236 ;
  assign n41302 = ~n41300 & ~n41301 ;
  assign n41282 = ~n41255 & n41256 ;
  assign n41271 = n40519 ^ n40518 ;
  assign n41272 = n41271 ^ n40116 ;
  assign n41273 = n41272 ^ n41243 ;
  assign n41274 = n41273 ^ n41271 ;
  assign n41275 = ~n41245 & ~n41274 ;
  assign n41276 = n41275 ^ n41272 ;
  assign n41277 = n41276 ^ n40463 ;
  assign n41278 = ~n39486 & ~n41277 ;
  assign n41279 = n41278 ^ n40463 ;
  assign n41266 = n41248 ^ n38764 ;
  assign n41267 = n41248 ^ n41239 ;
  assign n41268 = n41266 & ~n41267 ;
  assign n41269 = n41268 ^ n38764 ;
  assign n41270 = n41269 ^ n38956 ;
  assign n41280 = n41279 ^ n41270 ;
  assign n41262 = n41249 ^ x318 ;
  assign n41263 = ~n41254 & n41262 ;
  assign n41264 = n41263 ^ x318 ;
  assign n41265 = n41264 ^ x317 ;
  assign n41281 = n41280 ^ n41265 ;
  assign n41283 = n41282 ^ n41281 ;
  assign n41258 = n41257 ^ n41235 ;
  assign n41259 = ~n41236 & ~n41258 ;
  assign n41260 = n41259 ^ n40811 ;
  assign n41261 = n41260 ^ n40941 ;
  assign n41284 = n41283 ^ n41261 ;
  assign n41303 = n41302 ^ n41284 ;
  assign n41304 = n41301 ^ n41300 ;
  assign n41305 = n41299 ^ n41298 ;
  assign n41306 = n41297 ^ n41295 ;
  assign n41307 = n41294 ^ n41293 ;
  assign n41308 = n41292 ^ n41290 ;
  assign n41309 = n41289 ^ n41288 ;
  assign n41310 = n41287 ^ n41285 ;
  assign n41466 = ~n41284 & ~n41302 ;
  assign n41426 = n41283 ^ n41260 ;
  assign n41427 = n41283 ^ n40941 ;
  assign n41428 = n41426 & ~n41427 ;
  assign n41429 = n41428 ^ n40941 ;
  assign n41396 = ~n41281 & ~n41282 ;
  assign n41311 = n41280 ^ n41264 ;
  assign n41312 = n41280 ^ x317 ;
  assign n41313 = n41311 & ~n41312 ;
  assign n41314 = n41313 ^ x317 ;
  assign n41394 = n41314 ^ x316 ;
  assign n41325 = n40521 ^ n40520 ;
  assign n41321 = n40479 ^ n40463 ;
  assign n41320 = n41271 ^ n40479 ;
  assign n41322 = n41321 ^ n41320 ;
  assign n41323 = ~n41276 & ~n41322 ;
  assign n41324 = n41323 ^ n41321 ;
  assign n41326 = n41325 ^ n41324 ;
  assign n41327 = n39494 & ~n41326 ;
  assign n41328 = n41327 ^ n40479 ;
  assign n41315 = n41279 ^ n41269 ;
  assign n41316 = n41279 ^ n38956 ;
  assign n41317 = n41315 & ~n41316 ;
  assign n41318 = n41317 ^ n38956 ;
  assign n41319 = n41318 ^ n38969 ;
  assign n41329 = n41328 ^ n41319 ;
  assign n41395 = n41394 ^ n41329 ;
  assign n41424 = n41396 ^ n41395 ;
  assign n41425 = n41424 ^ n40979 ;
  assign n41467 = n41429 ^ n41425 ;
  assign n41468 = n41466 & n41467 ;
  assign n41397 = ~n41395 & ~n41396 ;
  assign n41330 = n41329 ^ n41314 ;
  assign n41341 = n40523 ^ n40522 ;
  assign n41337 = n40622 ^ n40479 ;
  assign n41336 = n41325 ^ n40622 ;
  assign n41338 = n41337 ^ n41336 ;
  assign n41339 = ~n41324 & n41338 ;
  assign n41340 = n41339 ^ n41337 ;
  assign n41342 = n41341 ^ n41340 ;
  assign n41343 = n39502 & n41342 ;
  assign n41344 = n41343 ^ n40622 ;
  assign n41331 = n41328 ^ n41318 ;
  assign n41332 = n41328 ^ n38969 ;
  assign n41333 = ~n41331 & n41332 ;
  assign n41334 = n41333 ^ n38969 ;
  assign n41335 = n41334 ^ n38982 ;
  assign n41345 = n41344 ^ n41335 ;
  assign n41346 = n41345 ^ x316 ;
  assign n41347 = n41346 ^ n41345 ;
  assign n41348 = n41347 ^ n41314 ;
  assign n41349 = ~n41330 & n41348 ;
  assign n41350 = n41349 ^ n41346 ;
  assign n41393 = n41350 ^ x315 ;
  assign n41433 = n41397 ^ n41393 ;
  assign n41469 = n41433 ^ n41006 ;
  assign n41430 = n41429 ^ n41424 ;
  assign n41431 = n41425 & ~n41430 ;
  assign n41432 = n41431 ^ n40979 ;
  assign n41470 = n41469 ^ n41432 ;
  assign n41471 = ~n41468 & n41470 ;
  assign n41434 = n41433 ^ n41432 ;
  assign n41398 = n41393 & ~n41397 ;
  assign n41358 = n41341 ^ n40622 ;
  assign n41359 = ~n41340 & n41358 ;
  assign n41360 = n41359 ^ n40622 ;
  assign n41356 = n40526 ^ n40524 ;
  assign n41357 = n41356 ^ n40641 ;
  assign n41361 = n41360 ^ n41357 ;
  assign n41362 = n39509 & n41361 ;
  assign n41363 = n41362 ^ n40641 ;
  assign n41351 = n41344 ^ n41334 ;
  assign n41352 = n41344 ^ n38982 ;
  assign n41353 = n41351 & n41352 ;
  assign n41354 = n41353 ^ n38982 ;
  assign n41355 = n41354 ^ n38995 ;
  assign n41364 = n41363 ^ n41355 ;
  assign n41366 = n41364 ^ x315 ;
  assign n41365 = n41364 ^ n41345 ;
  assign n41367 = n41366 ^ n41365 ;
  assign n41368 = ~n41350 & n41367 ;
  assign n41369 = n41368 ^ n41366 ;
  assign n41392 = n41369 ^ x314 ;
  assign n41422 = n41398 ^ n41392 ;
  assign n41435 = n41422 ^ n41006 ;
  assign n41436 = n41435 ^ n41432 ;
  assign n41437 = n41436 ^ n41422 ;
  assign n41438 = ~n41434 & ~n41437 ;
  assign n41439 = n41438 ^ n41435 ;
  assign n41472 = n41439 ^ n41033 ;
  assign n41473 = ~n41471 & n41472 ;
  assign n41381 = n40528 ^ n40527 ;
  assign n41375 = n41360 ^ n41356 ;
  assign n41376 = n40767 ^ n40641 ;
  assign n41377 = n41376 ^ n40767 ;
  assign n41378 = n41377 ^ n41356 ;
  assign n41379 = ~n41375 & ~n41378 ;
  assign n41380 = n41379 ^ n41376 ;
  assign n41382 = n41381 ^ n41380 ;
  assign n41383 = n39516 & ~n41382 ;
  assign n41384 = n41383 ^ n40767 ;
  assign n41370 = n41363 ^ n41354 ;
  assign n41371 = n41363 ^ n38995 ;
  assign n41372 = n41370 & ~n41371 ;
  assign n41373 = n41372 ^ n38995 ;
  assign n41374 = n41373 ^ n39009 ;
  assign n41385 = n41384 ^ n41374 ;
  assign n41387 = n41385 ^ x314 ;
  assign n41386 = n41385 ^ n41364 ;
  assign n41388 = n41387 ^ n41386 ;
  assign n41389 = ~n41369 & n41388 ;
  assign n41390 = n41389 ^ n41387 ;
  assign n41442 = n41390 ^ x313 ;
  assign n41399 = ~n41392 & ~n41398 ;
  assign n41443 = n41442 ^ n41399 ;
  assign n41474 = n41443 ^ n41088 ;
  assign n41423 = n41422 ^ n41033 ;
  assign n41440 = ~n41423 & n41439 ;
  assign n41441 = n41440 ^ n41033 ;
  assign n41475 = n41474 ^ n41441 ;
  assign n41476 = n41473 & ~n41475 ;
  assign n41444 = n41443 ^ n41441 ;
  assign n41414 = n40530 ^ n40529 ;
  assign n41415 = n41414 ^ n40802 ;
  assign n41416 = n41415 ^ n41381 ;
  assign n41412 = n41381 ^ n40767 ;
  assign n41413 = n41380 & ~n41412 ;
  assign n41417 = n41416 ^ n41413 ;
  assign n41418 = n39523 & ~n41417 ;
  assign n41408 = n39207 ^ n39009 ;
  assign n41409 = n41408 ^ n40802 ;
  assign n41410 = n41409 ^ x312 ;
  assign n41405 = n41384 ^ n41373 ;
  assign n41406 = n41384 ^ n39009 ;
  assign n41407 = ~n41405 & ~n41406 ;
  assign n41411 = n41410 ^ n41407 ;
  assign n41419 = n41418 ^ n41411 ;
  assign n41400 = n41399 ^ n41385 ;
  assign n41403 = ~n41390 & n41400 ;
  assign n41391 = n41390 ^ n41385 ;
  assign n41401 = n41400 ^ n41391 ;
  assign n41402 = x313 & n41401 ;
  assign n41404 = n41403 ^ n41402 ;
  assign n41420 = n41419 ^ n41404 ;
  assign n41445 = n41420 ^ n41088 ;
  assign n41446 = n41445 ^ n41441 ;
  assign n41447 = n41446 ^ n41420 ;
  assign n41448 = ~n41444 & n41447 ;
  assign n41449 = n41448 ^ n41445 ;
  assign n41477 = n41449 ^ n41084 ;
  assign n41478 = ~n41476 & ~n41477 ;
  assign n41479 = n41108 ^ n40900 ;
  assign n41421 = n41420 ^ n41084 ;
  assign n41450 = ~n41421 & ~n41449 ;
  assign n41451 = n41450 ^ n41084 ;
  assign n41480 = n41479 ^ n41451 ;
  assign n41481 = n41478 & ~n41480 ;
  assign n41458 = n40902 ^ n40900 ;
  assign n41452 = n41451 ^ n41108 ;
  assign n41453 = n41121 ^ n40900 ;
  assign n41454 = n41453 ^ n41121 ;
  assign n41455 = n41454 ^ n41451 ;
  assign n41456 = ~n41452 & n41455 ;
  assign n41457 = n41456 ^ n41453 ;
  assign n41482 = n41458 ^ n41457 ;
  assign n41483 = ~n41481 & n41482 ;
  assign n41464 = n40904 ^ n40903 ;
  assign n41460 = n41158 ^ n41121 ;
  assign n41459 = n41458 ^ n41158 ;
  assign n41461 = n41460 ^ n41459 ;
  assign n41462 = ~n41457 & n41461 ;
  assign n41463 = n41462 ^ n41460 ;
  assign n41465 = n41464 ^ n41463 ;
  assign n41484 = n41483 ^ n41465 ;
  assign n41485 = n41482 ^ n41481 ;
  assign n41486 = n41480 ^ n41478 ;
  assign n41487 = n41477 ^ n41476 ;
  assign n41488 = n41475 ^ n41473 ;
  assign n41489 = n41472 ^ n41471 ;
  assign n41490 = n41470 ^ n41468 ;
  assign n41491 = n41467 ^ n41466 ;
  assign n41497 = n41189 ^ n41158 ;
  assign n41496 = n41464 ^ n41189 ;
  assign n41498 = n41497 ^ n41496 ;
  assign n41499 = n41463 & n41498 ;
  assign n41500 = n41499 ^ n41497 ;
  assign n41504 = n40908 ^ n40907 ;
  assign n41506 = n41504 ^ n41189 ;
  assign n41501 = n40906 ^ n40905 ;
  assign n41505 = n41504 ^ n41501 ;
  assign n41507 = n41506 ^ n41505 ;
  assign n41508 = n41500 & ~n41507 ;
  assign n41509 = n41508 ^ n41506 ;
  assign n41513 = n41504 ^ n41246 ;
  assign n41514 = ~n41509 & ~n41513 ;
  assign n41515 = n41514 ^ n41246 ;
  assign n41512 = n40911 ^ n40909 ;
  assign n41516 = n41515 ^ n41512 ;
  assign n41520 = n41326 ^ n41277 ;
  assign n41519 = n41515 ^ n41326 ;
  assign n41521 = n41520 ^ n41519 ;
  assign n41522 = ~n41516 & ~n41521 ;
  assign n41523 = n41522 ^ n41520 ;
  assign n41528 = n41342 ^ n41326 ;
  assign n41524 = n40913 ^ n40912 ;
  assign n41527 = n41524 ^ n41342 ;
  assign n41529 = n41528 ^ n41527 ;
  assign n41530 = n41523 & ~n41529 ;
  assign n41531 = n41530 ^ n41528 ;
  assign n41532 = n40916 ^ n40914 ;
  assign n41537 = n41532 ^ n41342 ;
  assign n41538 = ~n41531 & ~n41537 ;
  assign n41539 = n41538 ^ n41342 ;
  assign n41535 = n40918 ^ n40917 ;
  assign n41543 = n41539 ^ n41535 ;
  assign n41544 = n41382 ^ n41361 ;
  assign n41545 = n41544 ^ n41382 ;
  assign n41546 = n41545 ^ n41535 ;
  assign n41547 = ~n41543 & n41546 ;
  assign n41548 = n41547 ^ n41544 ;
  assign n41551 = n41382 & n41548 ;
  assign n41495 = ~n41465 & n41483 ;
  assign n41502 = n41501 ^ n41500 ;
  assign n41503 = n41495 & n41502 ;
  assign n41510 = n41509 ^ n41246 ;
  assign n41511 = n41503 & n41510 ;
  assign n41517 = n41516 ^ n41277 ;
  assign n41518 = n41511 & ~n41517 ;
  assign n41525 = n41524 ^ n41523 ;
  assign n41526 = n41518 & n41525 ;
  assign n41533 = n41532 ^ n41531 ;
  assign n41534 = ~n41526 & ~n41533 ;
  assign n41536 = n41535 ^ n41361 ;
  assign n41540 = n41539 ^ n41536 ;
  assign n41541 = ~n41534 & n41540 ;
  assign n41494 = n40921 ^ n40919 ;
  assign n41542 = n41541 ^ n41494 ;
  assign n41549 = n41548 ^ n41494 ;
  assign n41550 = n41542 & n41549 ;
  assign n41552 = n41551 ^ n41550 ;
  assign n41492 = n40923 ^ n40922 ;
  assign n41493 = n41492 ^ n41417 ;
  assign n41553 = n41552 ^ n41493 ;
  assign n41554 = n41549 ^ n41541 ;
  assign n41555 = n41540 ^ n41534 ;
  assign n41556 = n41533 ^ n41526 ;
  assign n41557 = n41525 ^ n41518 ;
  assign n41558 = n41517 ^ n41511 ;
  assign n41559 = n41510 ^ n41503 ;
  assign n41560 = n41502 ^ n41495 ;
  assign n41561 = ~n40684 & n40692 ;
  assign n41562 = n40704 & n41561 ;
  assign n41563 = ~n40710 & n41562 ;
  assign n41564 = ~n40714 & n41563 ;
  assign n41565 = n40679 & n41564 ;
  assign n41566 = n41565 ^ n40675 ;
  assign n41567 = n41564 ^ n40679 ;
  assign n41568 = n41563 ^ n40714 ;
  assign n41569 = n41562 ^ n40710 ;
  assign n41570 = n41561 ^ n40704 ;
  assign n41571 = n40692 ^ n40684 ;
  assign n41572 = ~n40675 & n41565 ;
  assign n41573 = ~n40671 & ~n41572 ;
  assign n41574 = ~n40666 & n41573 ;
  assign n41575 = ~n40662 & ~n41574 ;
  assign n41576 = ~n40743 & n41575 ;
  assign n41577 = ~n40658 & n41576 ;
  assign n41578 = n40779 & ~n41577 ;
  assign n41579 = n40811 & ~n41578 ;
  assign n41580 = n41579 ^ n40941 ;
  assign n41581 = n41578 ^ n40811 ;
  assign n41582 = n41577 ^ n40779 ;
  assign n41583 = n41576 ^ n40658 ;
  assign n41584 = n41575 ^ n40743 ;
  assign n41585 = n41574 ^ n40662 ;
  assign n41586 = n41573 ^ n40666 ;
  assign n41587 = n41572 ^ n40671 ;
  assign n41588 = n40941 & n41579 ;
  assign n41589 = ~n40979 & ~n41588 ;
  assign n41590 = ~n41006 & ~n41589 ;
  assign n41591 = n41033 & ~n41590 ;
  assign n41592 = ~n41088 & ~n41591 ;
  assign n41593 = n41084 & n41592 ;
  assign n41594 = n41108 & n41593 ;
  assign n41595 = n41121 & ~n41594 ;
  assign n41596 = n41595 ^ n41158 ;
  assign n41597 = n41594 ^ n41121 ;
  assign n41598 = n41593 ^ n41108 ;
  assign n41599 = n41592 ^ n41084 ;
  assign n41600 = n41591 ^ n41088 ;
  assign n41601 = n41590 ^ n41033 ;
  assign n41602 = n41589 ^ n41006 ;
  assign n41603 = n41588 ^ n40979 ;
  assign n41604 = ~n41158 & ~n41595 ;
  assign n41605 = n41189 & ~n41604 ;
  assign n41606 = ~n41246 & n41605 ;
  assign n41607 = n41277 & n41606 ;
  assign n41608 = ~n41326 & ~n41607 ;
  assign n41609 = n41342 & n41608 ;
  assign n41610 = ~n41361 & ~n41609 ;
  assign n41611 = n41382 & n41610 ;
  assign n41612 = n41611 ^ n41417 ;
  assign n41613 = n41610 ^ n41382 ;
  assign n41614 = n41609 ^ n41361 ;
  assign n41615 = n41608 ^ n41342 ;
  assign n41616 = n41607 ^ n41326 ;
  assign n41617 = n41606 ^ n41277 ;
  assign n41618 = n41605 ^ n41246 ;
  assign n41619 = n41604 ^ n41189 ;
  assign n41620 = ~n40202 & ~n40209 ;
  assign n41621 = ~n40215 & ~n41620 ;
  assign n41622 = ~n40191 & ~n41621 ;
  assign n41623 = ~n40227 & n41622 ;
  assign n41624 = ~n40187 & n41623 ;
  assign n41625 = n41624 ^ n40183 ;
  assign n41626 = n41623 ^ n40187 ;
  assign n41627 = n41622 ^ n40227 ;
  assign n41628 = n41621 ^ n40191 ;
  assign n41629 = n41620 ^ n40215 ;
  assign n41630 = n40209 ^ n40202 ;
  assign n41631 = ~n40183 & ~n41624 ;
  assign n41632 = ~n40178 & n41631 ;
  assign n41633 = n40174 & n41632 ;
  assign n41634 = n40245 & ~n41633 ;
  assign n41635 = ~n40169 & ~n41634 ;
  assign n41636 = ~n40165 & ~n41635 ;
  assign n41637 = n40161 & ~n41636 ;
  assign n41638 = ~n40157 & ~n41637 ;
  assign n41639 = n41638 ^ n40153 ;
  assign n41640 = n41637 ^ n40157 ;
  assign n41641 = n41636 ^ n40161 ;
  assign n41642 = n41635 ^ n40165 ;
  assign n41643 = n41634 ^ n40169 ;
  assign n41644 = n41633 ^ n40245 ;
  assign n41645 = n41632 ^ n40174 ;
  assign n41646 = n41631 ^ n40178 ;
  assign n41647 = ~n40153 & ~n41638 ;
  assign n41648 = ~n40148 & n41647 ;
  assign n41649 = n40144 & ~n41648 ;
  assign n41650 = n40139 & ~n41649 ;
  assign n41651 = n40135 & n41650 ;
  assign n41652 = n40280 & ~n41651 ;
  assign n41653 = ~n40131 & n41652 ;
  assign n41654 = ~n40127 & ~n41653 ;
  assign n41655 = n41654 ^ n40123 ;
  assign n41656 = n41653 ^ n40127 ;
  assign n41657 = n41652 ^ n40131 ;
  assign n41658 = n41651 ^ n40280 ;
  assign n41659 = n41650 ^ n40135 ;
  assign n41660 = n41649 ^ n40139 ;
  assign n41661 = n41648 ^ n40144 ;
  assign n41662 = n41647 ^ n40148 ;
  assign n41663 = ~n40123 & n41654 ;
  assign n41664 = n40119 & n41663 ;
  assign n41665 = ~n40116 & n41664 ;
  assign n41666 = n40463 & n41665 ;
  assign n41667 = ~n40479 & n41666 ;
  assign n41668 = ~n40622 & ~n41667 ;
  assign n41669 = ~n40641 & ~n41668 ;
  assign n41670 = n40767 & n41669 ;
  assign n41671 = n41670 ^ n40802 ;
  assign n41672 = n41669 ^ n40767 ;
  assign n41673 = n41668 ^ n40641 ;
  assign n41674 = n41667 ^ n40622 ;
  assign n41675 = n41666 ^ n40479 ;
  assign n41676 = n41665 ^ n40463 ;
  assign n41677 = n41664 ^ n40116 ;
  assign n41678 = n41663 ^ n40119 ;
  assign y0 = n39322 ;
  assign y1 = n39323 ;
  assign y2 = ~n39324 ;
  assign y3 = ~n39325 ;
  assign y4 = ~n39326 ;
  assign y5 = ~n39327 ;
  assign y6 = ~n39328 ;
  assign y7 = ~n39308 ;
  assign y8 = n39388 ;
  assign y9 = ~n39389 ;
  assign y10 = n39390 ;
  assign y11 = n39391 ;
  assign y12 = n39392 ;
  assign y13 = n39393 ;
  assign y14 = ~n39394 ;
  assign y15 = n39395 ;
  assign y16 = n39455 ;
  assign y17 = ~n39456 ;
  assign y18 = n39457 ;
  assign y19 = ~n39458 ;
  assign y20 = n39459 ;
  assign y21 = n39460 ;
  assign y22 = ~n39461 ;
  assign y23 = ~n39462 ;
  assign y24 = ~n39524 ;
  assign y25 = n39525 ;
  assign y26 = ~n39526 ;
  assign y27 = n39527 ;
  assign y28 = ~n39528 ;
  assign y29 = ~n39529 ;
  assign y30 = ~n39530 ;
  assign y31 = n39531 ;
  assign y32 = ~n41067 ;
  assign y33 = ~n41068 ;
  assign y34 = ~n41069 ;
  assign y35 = n41070 ;
  assign y36 = n41071 ;
  assign y37 = n41072 ;
  assign y38 = ~n41073 ;
  assign y39 = ~n41051 ;
  assign y40 = ~n41303 ;
  assign y41 = n41304 ;
  assign y42 = ~n41305 ;
  assign y43 = n41306 ;
  assign y44 = ~n41307 ;
  assign y45 = ~n41308 ;
  assign y46 = ~n41309 ;
  assign y47 = ~n41310 ;
  assign y48 = n41484 ;
  assign y49 = n41485 ;
  assign y50 = ~n41486 ;
  assign y51 = n41487 ;
  assign y52 = n41488 ;
  assign y53 = n41489 ;
  assign y54 = ~n41490 ;
  assign y55 = ~n41491 ;
  assign y56 = n41553 ;
  assign y57 = ~n41554 ;
  assign y58 = n41555 ;
  assign y59 = n41556 ;
  assign y60 = ~n41557 ;
  assign y61 = n41558 ;
  assign y62 = ~n41559 ;
  assign y63 = ~n41560 ;
  assign y64 = n41566 ;
  assign y65 = ~n41567 ;
  assign y66 = n41568 ;
  assign y67 = n41569 ;
  assign y68 = ~n41570 ;
  assign y69 = n41571 ;
  assign y70 = n40692 ;
  assign y71 = n40688 ;
  assign y72 = ~n41580 ;
  assign y73 = n41581 ;
  assign y74 = ~n41582 ;
  assign y75 = n41583 ;
  assign y76 = n41584 ;
  assign y77 = ~n41585 ;
  assign y78 = ~n41586 ;
  assign y79 = n41587 ;
  assign y80 = ~n41596 ;
  assign y81 = ~n41597 ;
  assign y82 = ~n41598 ;
  assign y83 = ~n41599 ;
  assign y84 = ~n41600 ;
  assign y85 = ~n41601 ;
  assign y86 = ~n41602 ;
  assign y87 = n41603 ;
  assign y88 = ~n41612 ;
  assign y89 = n41613 ;
  assign y90 = n41614 ;
  assign y91 = ~n41615 ;
  assign y92 = ~n41616 ;
  assign y93 = n41617 ;
  assign y94 = ~n41618 ;
  assign y95 = ~n41619 ;
  assign y96 = n41625 ;
  assign y97 = n41626 ;
  assign y98 = n41627 ;
  assign y99 = ~n41628 ;
  assign y100 = n41629 ;
  assign y101 = ~n41630 ;
  assign y102 = ~n40202 ;
  assign y103 = ~n40196 ;
  assign y104 = n41639 ;
  assign y105 = ~n41640 ;
  assign y106 = ~n41641 ;
  assign y107 = ~n41642 ;
  assign y108 = n41643 ;
  assign y109 = n41644 ;
  assign y110 = n41645 ;
  assign y111 = ~n41646 ;
  assign y112 = ~n41655 ;
  assign y113 = n41656 ;
  assign y114 = n41657 ;
  assign y115 = n41658 ;
  assign y116 = n41659 ;
  assign y117 = ~n41660 ;
  assign y118 = n41661 ;
  assign y119 = ~n41662 ;
  assign y120 = n41671 ;
  assign y121 = n41672 ;
  assign y122 = n41673 ;
  assign y123 = ~n41674 ;
  assign y124 = ~n41675 ;
  assign y125 = n41676 ;
  assign y126 = ~n41677 ;
  assign y127 = n41678 ;
endmodule
