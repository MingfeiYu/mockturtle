module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n197 , n198 , n199 , n200 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n265 , n266 , n267 , n268 , n269 ;
  assign n65 = x59 ^ x27 ;
  assign n69 = x27 & ~x59 ;
  assign n67 = x25 & x57 ;
  assign n66 = x58 ^ x57 ;
  assign n68 = n67 ^ n66 ;
  assign n70 = n69 ^ n68 ;
  assign n73 = x59 ^ x26 ;
  assign n71 = x59 ^ x57 ;
  assign n72 = n71 ^ n67 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~n70 & ~n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = ~n65 & n76 ;
  assign n78 = n77 ^ x27 ;
  assign n79 = x28 & ~x60 ;
  assign n80 = ~x31 & x63 ;
  assign n81 = ~n79 & n80 ;
  assign n82 = n81 ^ x29 ;
  assign n83 = n81 ^ n79 ;
  assign n84 = ~x61 & ~n83 ;
  assign n85 = n82 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = x30 & ~x62 ;
  assign n88 = ~n86 & n87 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = n78 & ~n89 ;
  assign n134 = n67 ^ x25 ;
  assign n135 = ~n69 & ~n134 ;
  assign n136 = x26 & ~x58 ;
  assign n137 = n135 & n136 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = ~x24 & n138 ;
  assign n91 = x20 & ~x52 ;
  assign n92 = x21 & ~x53 ;
  assign n94 = ~x22 & x54 ;
  assign n93 = x54 ^ x22 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = ~n92 & ~n95 ;
  assign n97 = x23 & ~x55 ;
  assign n98 = n96 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = ~n91 & n99 ;
  assign n102 = x16 & ~x48 ;
  assign n101 = x48 ^ x16 ;
  assign n103 = n102 ^ n101 ;
  assign n105 = x17 & ~x49 ;
  assign n104 = x49 ^ x17 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = ~n103 & ~n106 ;
  assign n109 = ~x18 & x50 ;
  assign n108 = x50 ^ x18 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = ~n105 & ~n110 ;
  assign n112 = x19 & ~x51 ;
  assign n113 = n111 & n112 ;
  assign n114 = n113 ^ n111 ;
  assign n115 = ~n107 & n114 ;
  assign n116 = x51 ^ x19 ;
  assign n117 = n109 ^ x51 ;
  assign n118 = ~n116 & n117 ;
  assign n119 = n118 ^ x51 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = n100 & ~n120 ;
  assign n122 = x52 ^ x20 ;
  assign n123 = n122 ^ n91 ;
  assign n124 = x53 ^ x21 ;
  assign n125 = n124 ^ n92 ;
  assign n126 = ~n123 & ~n125 ;
  assign n127 = n99 & ~n126 ;
  assign n128 = x55 ^ x23 ;
  assign n129 = n94 ^ x55 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = n130 ^ x55 ;
  assign n132 = ~n127 & ~n131 ;
  assign n133 = ~n121 & n132 ;
  assign n140 = n139 ^ n133 ;
  assign n141 = x56 & n138 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = ~n140 & n142 ;
  assign n144 = n143 ^ n139 ;
  assign n145 = n90 & ~n144 ;
  assign n146 = n145 ^ n89 ;
  assign n147 = x63 ^ x31 ;
  assign n149 = x60 ^ x28 ;
  assign n150 = n149 ^ n79 ;
  assign n151 = n150 ^ x62 ;
  assign n148 = x62 ^ x29 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = x62 ^ x61 ;
  assign n154 = n153 ^ n151 ;
  assign n155 = ~n152 & n154 ;
  assign n156 = n155 ^ n151 ;
  assign n158 = x63 ^ x30 ;
  assign n157 = x63 ^ x62 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = ~n147 & ~n161 ;
  assign n163 = n162 ^ x31 ;
  assign n164 = x47 ^ x15 ;
  assign n166 = x14 & ~x46 ;
  assign n165 = x46 ^ x14 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = n167 ^ x47 ;
  assign n169 = ~n164 & ~n168 ;
  assign n170 = n169 ^ x15 ;
  assign n171 = x45 ^ x13 ;
  assign n173 = x12 & ~x44 ;
  assign n172 = x44 ^ x12 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = n174 ^ x45 ;
  assign n176 = ~n171 & ~n175 ;
  assign n177 = n176 ^ x13 ;
  assign n178 = ~n171 & ~n173 ;
  assign n179 = ~n164 & ~n166 ;
  assign n180 = x42 ^ x10 ;
  assign n181 = x43 ^ x11 ;
  assign n182 = ~n180 & ~n181 ;
  assign n184 = ~x9 & x41 ;
  assign n183 = x41 ^ x9 ;
  assign n185 = n184 ^ n183 ;
  assign n188 = ~x8 & ~n185 ;
  assign n189 = n182 & n188 ;
  assign n186 = x40 & ~n185 ;
  assign n187 = n182 & n186 ;
  assign n190 = n189 ^ n187 ;
  assign n229 = n187 ^ x39 ;
  assign n191 = x38 ^ x6 ;
  assign n192 = x5 & x37 ;
  assign n193 = n192 ^ x5 ;
  assign n194 = x36 ^ x4 ;
  assign n197 = x34 ^ x2 ;
  assign n199 = x34 ^ x1 ;
  assign n198 = x34 ^ x33 ;
  assign n200 = n199 ^ n198 ;
  assign n202 = x0 & ~x32 ;
  assign n203 = n202 ^ x1 ;
  assign n204 = ~n200 & n203 ;
  assign n205 = n204 ^ n199 ;
  assign n206 = ~n197 & n205 ;
  assign n195 = x35 ^ x2 ;
  assign n207 = n206 ^ n195 ;
  assign n209 = x36 ^ x3 ;
  assign n208 = x36 ^ x35 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n207 & ~n210 ;
  assign n212 = n211 ^ n209 ;
  assign n213 = ~n194 & n212 ;
  assign n214 = n213 ^ x4 ;
  assign n215 = ~n193 & ~n214 ;
  assign n216 = ~n191 & n215 ;
  assign n221 = x7 & ~x39 ;
  assign n222 = n221 ^ n191 ;
  assign n223 = n192 ^ x37 ;
  assign n224 = n223 ^ x6 ;
  assign n225 = ~n222 & ~n224 ;
  assign n226 = n225 ^ x6 ;
  assign n227 = ~n216 & n226 ;
  assign n228 = n227 ^ n187 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n187 ^ x7 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = ~n230 & ~n232 ;
  assign n234 = n233 ^ n229 ;
  assign n235 = n190 & ~n234 ;
  assign n236 = n235 ^ n189 ;
  assign n240 = n184 ^ x43 ;
  assign n237 = x43 ^ x42 ;
  assign n241 = n240 ^ n237 ;
  assign n242 = ~n180 & n241 ;
  assign n243 = n242 ^ n237 ;
  assign n244 = ~n181 & n243 ;
  assign n245 = n244 ^ x43 ;
  assign n246 = ~n236 & ~n245 ;
  assign n247 = n179 & ~n246 ;
  assign n248 = n178 & n247 ;
  assign n249 = n248 ^ n179 ;
  assign n250 = n177 & n249 ;
  assign n251 = n250 ^ n179 ;
  assign n252 = n170 & ~n251 ;
  assign n253 = ~n102 & ~n252 ;
  assign n254 = n114 & n253 ;
  assign n255 = n100 & n254 ;
  assign n256 = ~n89 & n255 ;
  assign n257 = ~n163 & n256 ;
  assign n265 = ~n141 & n257 ;
  assign n266 = ~n139 & n265 ;
  assign n267 = n266 ^ n139 ;
  assign n258 = n257 ^ n163 ;
  assign n259 = n258 ^ n139 ;
  assign n268 = n267 ^ n259 ;
  assign n269 = n146 & ~n268 ;
  assign y0 = ~n269 ;
endmodule
