module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n95 , n96 , n97 , n100 , n101 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n117 , n124 , n125 , n126 , n131 , n132 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n150 , n151 , n152 , n155 , n156 , n157 , n158 , n159 , n162 , n163 , n164 , n165 , n167 , n168 , n169 , n172 , n173 , n176 , n178 , n179 , n181 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n207 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 ;
  assign n35 = x5 ^ x3 ;
  assign n28 = x1 & x4 ;
  assign n26 = x3 ^ x2 ;
  assign n24 = x3 ^ x1 ;
  assign n25 = n24 ^ x0 ;
  assign n27 = n26 ^ n25 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~x5 & n29 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = ~x6 & n31 ;
  assign n23 = x4 ^ x2 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = ~x7 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = ~x8 & n36 ;
  assign n22 = x6 ^ x4 ;
  assign n38 = n37 ^ n22 ;
  assign n39 = ~x9 & n38 ;
  assign n20 = x6 ^ x5 ;
  assign n13 = x6 & x7 ;
  assign n15 = ~x8 & ~n13 ;
  assign n14 = n13 ^ x8 ;
  assign n16 = n15 ^ n14 ;
  assign n18 = ~x9 & ~n16 ;
  assign n12 = x7 ^ x6 ;
  assign n17 = n16 ^ n12 ;
  assign n19 = n18 ^ n17 ;
  assign n21 = n20 ^ n19 ;
  assign n40 = n39 ^ n21 ;
  assign n41 = ~x10 & ~n40 ;
  assign n42 = n41 ^ n19 ;
  assign n43 = ~x7 & ~x8 ;
  assign n58 = ~x2 & ~x3 ;
  assign n59 = n58 ^ n26 ;
  assign n53 = x1 & x2 ;
  assign n46 = ~x0 & n28 ;
  assign n44 = x2 & x4 ;
  assign n45 = n44 ^ x1 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n47 ^ x3 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = x5 & n54 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = n56 ^ x4 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n60 ^ n56 ;
  assign n64 = ~x9 & n61 ;
  assign n65 = n64 ^ n56 ;
  assign n66 = x6 & ~n65 ;
  assign n67 = n66 ^ n56 ;
  assign n68 = n43 & ~n67 ;
  assign n81 = ~x5 & ~x6 ;
  assign n82 = n81 ^ n20 ;
  assign n83 = n82 ^ x7 ;
  assign n70 = x4 & x5 ;
  assign n71 = n70 ^ x6 ;
  assign n84 = n83 ^ n71 ;
  assign n69 = x9 ^ x8 ;
  assign n73 = x3 & x4 ;
  assign n72 = n71 ^ x5 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n71 ;
  assign n78 = x7 & ~n75 ;
  assign n79 = n78 ^ n71 ;
  assign n80 = ~n69 & ~n79 ;
  assign n85 = n84 ^ n80 ;
  assign n86 = ~x9 & ~n85 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = ~x10 & ~n87 ;
  assign n89 = ~n68 & n88 ;
  assign n90 = x10 & ~n15 ;
  assign n91 = ~n18 & n90 ;
  assign n92 = ~n89 & ~n91 ;
  assign n217 = x5 & n13 ;
  assign n216 = n16 ^ x8 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = ~x10 & n218 ;
  assign n220 = n219 ^ n16 ;
  assign n106 = x8 & ~n12 ;
  assign n93 = x8 ^ x7 ;
  assign n95 = n93 ^ n70 ;
  assign n96 = n95 ^ x3 ;
  assign n117 = x6 ^ x3 ;
  assign n97 = n95 ^ n71 ;
  assign n100 = n117 ^ n97 ;
  assign n101 = n96 & ~n100 ;
  assign n107 = n106 ^ n101 ;
  assign n108 = n107 ^ n97 ;
  assign n109 = n106 ^ x6 ;
  assign n110 = n109 ^ n97 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = n71 & n111 ;
  assign n113 = n112 ^ n106 ;
  assign n114 = n113 ^ x8 ;
  assign n139 = n13 ^ x3 ;
  assign n185 = ~n13 & ~n139 ;
  assign n141 = x6 & n70 ;
  assign n142 = ~n59 & n141 ;
  assign n143 = ~x7 & ~n142 ;
  assign n144 = n143 ^ n13 ;
  assign n145 = n144 ^ n139 ;
  assign n140 = n139 ^ x5 ;
  assign n146 = n145 ^ n140 ;
  assign n124 = x6 ^ x2 ;
  assign n131 = x4 & n124 ;
  assign n125 = n124 ^ n20 ;
  assign n126 = n125 ^ n22 ;
  assign n132 = n131 ^ n126 ;
  assign n135 = n131 ^ x4 ;
  assign n136 = ~n117 & n135 ;
  assign n137 = n136 ^ x6 ;
  assign n138 = n132 & ~n137 ;
  assign n147 = n146 ^ n138 ;
  assign n172 = n147 ^ n143 ;
  assign n173 = n172 ^ n139 ;
  assign n186 = n185 ^ n173 ;
  assign n148 = n147 ^ n139 ;
  assign n187 = n186 ^ n148 ;
  assign n188 = n187 ^ x3 ;
  assign n150 = x3 & ~x6 ;
  assign n151 = n44 & n150 ;
  assign n167 = n151 ^ n144 ;
  assign n155 = x3 & ~x5 ;
  assign n156 = n155 ^ x6 ;
  assign n157 = x4 & ~n156 ;
  assign n152 = n151 ^ n20 ;
  assign n158 = n157 ^ n152 ;
  assign n159 = x3 ^ x0 ;
  assign n162 = x5 & n159 ;
  assign n163 = n162 ^ x0 ;
  assign n164 = x1 & n163 ;
  assign n165 = n158 & ~n164 ;
  assign n168 = n167 ^ n165 ;
  assign n203 = n168 ^ n139 ;
  assign n181 = n203 ^ n173 ;
  assign n189 = n181 ^ n148 ;
  assign n190 = n189 ^ x3 ;
  assign n191 = ~n188 & ~n190 ;
  assign n204 = n203 ^ n147 ;
  assign n205 = n204 ^ n144 ;
  assign n207 = n205 ^ n13 ;
  assign n176 = n207 ^ n148 ;
  assign n192 = n203 ^ n176 ;
  assign n178 = n176 ^ x3 ;
  assign n193 = n192 ^ n178 ;
  assign n195 = n204 ^ n178 ;
  assign n196 = n193 & n195 ;
  assign n197 = n191 & n196 ;
  assign n198 = n197 ^ n185 ;
  assign n199 = n198 ^ n181 ;
  assign n179 = n207 ^ n178 ;
  assign n200 = n199 ^ n179 ;
  assign n169 = n168 ^ n147 ;
  assign n201 = n200 ^ n169 ;
  assign n202 = n201 ^ n178 ;
  assign n209 = n202 ^ n143 ;
  assign n210 = n209 ^ x3 ;
  assign n211 = n210 ^ n207 ;
  assign n212 = ~x8 & ~n211 ;
  assign n213 = ~n114 & n212 ;
  assign n214 = n213 ^ n114 ;
  assign n215 = ~x10 & n214 ;
  assign n221 = n220 ^ n215 ;
  assign n222 = n220 ^ x9 ;
  assign n223 = n222 ^ x10 ;
  assign n224 = n223 ^ n215 ;
  assign n225 = ~n221 & ~n224 ;
  assign n226 = n225 ^ n222 ;
  assign n227 = ~x9 & ~x10 ;
  assign n228 = ~x3 & n227 ;
  assign n232 = ~x2 & ~n16 ;
  assign n233 = n70 & n232 ;
  assign n229 = x4 & n81 ;
  assign n230 = n229 ^ n81 ;
  assign n231 = n43 & n230 ;
  assign n234 = n233 ^ n231 ;
  assign n235 = n228 & n234 ;
  assign n236 = ~n69 & n217 ;
  assign n237 = ~x10 & n236 ;
  assign n240 = n237 ^ x10 ;
  assign n238 = ~x8 & ~n73 ;
  assign n239 = n237 & n238 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = ~x9 & ~n241 ;
  assign n243 = ~n58 & n70 ;
  assign n244 = n13 & n243 ;
  assign n246 = n229 ^ x6 ;
  assign n245 = n151 & n164 ;
  assign n247 = n246 ^ n245 ;
  assign n254 = n43 & ~n142 ;
  assign n249 = n247 & n254 ;
  assign n250 = n249 ^ x8 ;
  assign n251 = ~n244 & n250 ;
  assign n252 = n242 & n251 ;
  assign n253 = n252 ^ n241 ;
  assign n255 = n227 & n254 ;
  assign n257 = n81 & ~n245 ;
  assign n258 = n255 & n257 ;
  assign n256 = n255 ^ n227 ;
  assign n259 = n258 ^ n256 ;
  assign n260 = x8 & n244 ;
  assign n261 = n259 & n260 ;
  assign n262 = n261 ^ n259 ;
  assign y0 = ~n42 ;
  assign y1 = ~n92 ;
  assign y2 = ~n226 ;
  assign y3 = ~n235 ;
  assign y4 = n253 ;
  assign y5 = ~n262 ;
  assign y6 = ~n255 ;
endmodule
