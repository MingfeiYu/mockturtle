module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1357 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1373 , n1374 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1404 , n1405 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1482 , n1483 , n1484 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1540 , n1541 , n1545 , n1546 , n1547 , n1548 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1649 , n1650 , n1651 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1816 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1869 , n1870 , n1871 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1885 , n1886 , n1887 , n1888 , n1889 , n1892 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2094 , n2095 , n2101 , n2102 , n2103 , n2104 , n2105 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2118 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2165 , n2166 , n2169 , n2170 , n2171 , n2172 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2233 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2301 , n2302 , n2303 , n2304 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2314 , n2317 , n2318 , n2319 , n2320 , n2321 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2346 , n2347 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2396 , n2397 , n2398 , n2399 , n2401 , n2402 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2453 , n2454 , n2455 , n2456 , n2458 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2492 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2767 , n2769 , n2770 , n2771 , n2772 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2830 , n2832 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2916 , n2917 , n2918 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2939 , n2940 , n2941 , n2943 , n2944 , n2945 , n2947 , n2948 , n2949 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2968 , n2969 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3236 , n3237 , n3238 , n3239 , n3240 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3270 , n3271 , n3272 , n3273 , n3274 , n3276 , n3277 , n3278 , n3279 , n3280 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3311 , n3312 , n3317 , n3318 , n3319 , n3320 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3376 , n3385 , n3394 , n3395 , n3396 , n3397 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3429 , n3430 , n3431 , n3433 , n3434 , n3435 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3459 , n3462 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3474 , n3477 , n3478 , n3479 , n3480 , n3481 , n3483 , n3484 , n3485 , n3486 , n3490 , n3491 , n3492 , n3493 , n3494 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3521 , n3522 , n3523 , n3524 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3557 , n3560 , n3561 , n3562 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3600 , n3601 , n3602 , n3603 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3643 , n3644 , n3645 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3687 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3748 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3835 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3869 , n3870 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4011 , n4012 , n4013 , n4014 , n4019 , n4020 , n4021 , n4022 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4082 , n4083 , n4084 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4103 , n4104 , n4109 , n4110 , n4111 , n4112 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4144 , n4145 , n4146 , n4147 , n4148 , n4150 , n4159 , n4168 , n4169 , n4170 , n4171 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4195 , n4196 , n4197 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4223 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4270 , n4271 , n4272 , n4274 , n4275 , n4276 , n4277 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4386 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4413 , n4414 , n4415 , n4416 , n4417 , n4419 , n4420 , n4421 , n4423 , n4424 , n4425 , n4426 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4488 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4525 , n4526 , n4527 , n4528 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4687 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4699 , n4701 , n4710 , n4719 , n4720 , n4721 , n4722 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4746 , n4747 , n4748 , n4751 , n4752 , n4753 , n4755 , n4756 , n4757 , n4766 , n4775 , n4776 , n4777 , n4778 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4802 , n4803 , n4804 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4822 , n4823 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4905 , n4906 , n4907 , n4912 , n4913 , n4914 , n4915 , n4916 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5019 , n5020 , n5021 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5037 , n5038 , n5039 , n5040 , n5042 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5117 , n5118 , n5119 , n5120 , n5121 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5196 , n5197 , n5198 , n5199 , n5200 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5277 , n5278 , n5279 , n5284 , n5285 , n5286 , n5287 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5354 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5395 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5425 , n5430 , n5431 , n5432 , n5433 , n5434 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5460 , n5461 , n5462 , n5463 , n5464 , n5467 , n5468 , n5469 , n5470 , n5474 , n5475 , n5476 , n5477 , n5478 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5573 , n5576 , n5577 , n5578 , n5579 , n5580 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5632 , n5633 , n5634 , n5635 , n5636 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5670 , n5671 , n5672 , n5689 , n5690 , n5691 , n5692 , n5695 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5710 , n5711 , n5712 , n5726 , n5727 , n5728 , n5730 , n5731 , n5732 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5744 , n5745 , n5746 , n5747 , n5748 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5947 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5956 , n5959 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5968 , n5969 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6004 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6013 , n6016 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6025 , n6028 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6037 , n6038 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6051 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6060 , n6061 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6132 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6421 , n6422 , n6423 , n6424 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6622 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6632 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6756 , n6757 , n6758 , n6759 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6797 , n6798 , n6799 , n6800 , n6801 , n6803 , n6808 , n6809 , n6810 , n6811 , n6816 , n6830 , n6831 , n6832 , n6838 , n6839 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6860 , n6861 , n6862 , n6864 , n6865 , n6866 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6912 , n6913 , n6914 , n6915 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6928 , n6929 , n6930 , n6931 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7027 , n7028 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7049 , n7050 , n7051 , n7052 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7063 , n7064 , n7065 , n7066 , n7067 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7078 , n7079 , n7080 , n7081 , n7082 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7139 , n7140 , n7141 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7189 , n7190 , n7191 , n7194 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7219 , n7220 , n7221 , n7222 , n7223 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7237 , n7238 , n7239 , n7240 , n7242 , n7243 , n7246 , n7249 , n7250 , n7251 , n7252 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7264 , n7267 , n7268 , n7269 , n7270 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7284 , n7285 , n7286 , n7287 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7340 , n7343 , n7344 , n7345 , n7346 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7358 , n7361 , n7362 , n7363 , n7364 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7385 , n7388 , n7389 , n7390 , n7391 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7733 , n7736 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7796 , n7797 , n7799 , n7800 , n7805 , n7806 , n7807 , n7808 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8803 , n8804 , n8805 , n8806 , n8809 , n8810 , n8811 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8945 , n8946 , n8947 , n8948 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9010 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9035 , n9036 , n9037 , n9038 , n9041 , n9042 , n9043 , n9044 , n9047 , n9048 , n9049 , n9050 , n9053 , n9054 , n9055 , n9056 , n9059 , n9060 , n9061 , n9062 , n9065 , n9066 , n9067 , n9068 , n9071 , n9072 , n9073 , n9074 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9110 , n9111 , n9112 , n9113 , n9116 , n9117 , n9118 , n9119 , n9122 , n9123 , n9124 , n9125 , n9128 , n9129 , n9130 , n9131 , n9134 , n9135 , n9136 , n9137 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9166 , n9167 , n9168 , n9169 , n9172 , n9173 , n9174 , n9175 , n9178 , n9179 , n9180 , n9181 , n9184 , n9185 , n9186 , n9187 , n9190 , n9191 , n9192 , n9193 , n9196 , n9197 , n9198 , n9199 , n9202 , n9203 , n9204 , n9205 , n9208 , n9209 , n9210 , n9211 , n9214 , n9215 , n9216 , n9217 , n9220 , n9221 , n9222 , n9223 , n9226 , n9227 , n9228 , n9229 , n9232 , n9233 , n9234 , n9235 , n9238 , n9239 , n9240 , n9241 , n9244 , n9245 , n9246 , n9247 , n9250 , n9251 , n9252 , n9253 , n9256 , n9257 , n9258 , n9259 , n9262 , n9263 , n9264 , n9265 , n9268 , n9269 , n9270 , n9271 , n9274 , n9275 , n9276 , n9277 , n9280 , n9281 , n9282 , n9283 , n9286 , n9287 , n9288 , n9289 , n9292 , n9293 , n9294 , n9295 , n9298 , n9299 , n9300 , n9301 , n9304 , n9305 , n9306 , n9307 , n9310 , n9311 , n9312 , n9313 , n9316 , n9317 , n9318 , n9319 , n9322 , n9323 , n9324 , n9325 , n9328 , n9329 , n9330 , n9331 , n9334 , n9335 , n9336 , n9337 , n9340 , n9341 , n9342 , n9343 , n9346 , n9347 , n9348 , n9349 , n9352 , n9353 , n9354 , n9355 , n9358 , n9359 , n9360 , n9361 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9380 , n9381 , n9382 , n9383 , n9386 , n9387 , n9388 , n9389 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9484 , n9485 , n9486 , n9487 , n9488 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9538 , n9539 , n9540 , n9541 , n9542 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9562 , n9563 , n9564 , n9565 , n9566 , n9568 , n9570 , n9571 , n9573 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9612 , n9613 , n9614 , n9615 , n9616 , n9618 , n9620 , n9621 , n9623 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9672 , n9673 , n9674 , n9675 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9757 , n9758 , n9759 , n9760 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9772 , n9773 , n9774 , n9775 , n9776 , n9778 , n9780 , n9781 , n9783 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9846 , n9847 , n9848 , n9849 , n9850 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9870 , n9871 , n9872 , n9873 , n9874 , n9876 , n9878 , n9879 , n9880 , n9881 , n9882 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9944 , n9945 , n9946 , n9947 , n9948 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9968 , n9969 , n9970 , n9971 , n9972 , n9974 , n9976 , n9977 , n9979 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10022 , n10023 , n10024 , n10025 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10036 , n10037 , n10038 , n10039 , n10040 , n10042 , n10044 , n10045 , n10046 , n10047 , n10048 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10065 , n10066 , n10067 , n10068 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10171 , n10172 , n10173 , n10174 , n10177 , n10178 , n10179 , n10180 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10210 , n10211 , n10212 , n10213 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10225 , n10226 , n10227 , n10228 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10277 , n10278 , n10279 , n10280 , n10283 , n10284 , n10285 , n10286 , n10289 , n10290 , n10291 , n10292 , n10295 , n10296 , n10297 , n10298 , n10299 , n10301 , n10303 , n10304 , n10305 , n10306 , n10307 , n10310 , n10311 , n10312 , n10313 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10341 , n10342 , n10343 , n10344 , n10347 , n10348 , n10349 , n10350 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10398 , n10399 , n10400 , n10401 , n10404 , n10405 , n10406 , n10407 , n10410 , n10411 , n10412 , n10413 , n10416 , n10417 , n10418 , n10419 , n10422 , n10423 , n10424 , n10425 , n10428 , n10429 , n10430 , n10431 , n10434 , n10435 , n10436 , n10437 , n10440 , n10441 , n10442 , n10443 , n10446 , n10447 , n10448 , n10449 , n10452 , n10453 , n10454 , n10455 , n10458 , n10459 , n10460 , n10461 , n10464 , n10465 , n10466 , n10467 , n10470 , n10471 , n10472 , n10473 , n10476 , n10477 , n10478 , n10479 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10490 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10513 , n10514 , n10515 , n10516 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10532 , n10533 , n10534 , n10535 , n10538 , n10539 , n10540 , n10541 , n10542 , n10544 , n10548 , n10549 , n10550 , n10551 , n10554 , n10555 , n10556 , n10557 , n10558 , n10560 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10574 , n10575 , n10576 , n10577 , n10580 , n10581 , n10582 , n10583 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10594 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10617 , n10618 , n10619 , n10620 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10640 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10663 , n10664 , n10665 , n10666 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10686 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10709 , n10710 , n10711 , n10712 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10724 , n10725 , n10726 , n10727 , n10728 , n10730 , n10732 , n10733 , n10734 , n10735 , n10736 , n10739 , n10740 , n10741 , n10742 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10781 , n10782 , n10783 , n10784 , n10787 , n10788 , n10789 , n10790 , n10791 , n10793 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10829 , n10830 , n10831 , n10832 , n10833 , n10835 , n10837 , n10838 , n10839 , n10840 , n10841 , n10844 , n10845 , n10846 , n10847 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10878 , n10879 , n10880 , n10881 , n10882 , n10884 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10902 , n10903 , n10904 , n10905 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10917 , n10918 , n10919 , n10920 , n10921 , n10923 , n10925 , n10926 , n10927 , n10928 , n10929 , n10932 , n10933 , n10934 , n10935 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10963 , n10964 , n10965 , n10966 , n10967 , n10969 , n10971 , n10972 , n10973 , n10974 , n10975 , n10978 , n10979 , n10980 , n10981 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11031 , n11032 , n11033 , n11034 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11083 , n11084 , n11085 , n11086 , n11089 , n11090 , n11091 , n11092 , n11095 , n11096 , n11097 , n11098 , n11101 , n11102 , n11103 , n11104 , n11107 , n11108 , n11109 , n11110 , n11113 , n11114 , n11115 , n11116 , n11119 , n11120 , n11121 , n11122 , n11125 , n11126 , n11127 , n11128 , n11133 , n11134 , n11135 , n11136 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11149 , n11150 , n11151 , n11152 , n11155 , n11156 , n11157 , n11158 , n11159 , n11161 , n11165 , n11166 , n11167 , n11168 , n11171 , n11172 , n11173 , n11174 , n11175 , n11177 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11191 , n11192 , n11193 , n11194 , n11197 , n11198 , n11199 , n11200 , n11203 , n11204 , n11205 , n11206 , n11209 , n11210 , n11211 , n11212 , n11215 , n11216 , n11217 , n11218 , n11221 , n11222 , n11223 , n11224 , n11227 , n11228 , n11229 , n11230 , n11233 , n11234 , n11235 , n11236 , n11239 , n11240 , n11241 , n11242 , n11245 , n11246 , n11247 , n11248 , n11251 , n11252 , n11253 , n11254 , n11257 , n11258 , n11259 , n11264 , n11265 , n11266 , n11267 , n11270 , n11271 , n11272 , n11273 , n11276 , n11277 , n11278 , n11279 , n11282 , n11283 , n11284 , n11285 , n11288 , n11289 , n11290 , n11291 , n11294 , n11295 , n11296 , n11297 , n11300 , n11301 , n11302 , n11303 , n11306 , n11307 , n11308 , n11309 , n11312 , n11313 , n11314 , n11315 , n11318 , n11319 , n11320 , n11321 , n11324 , n11325 , n11326 , n11327 , n11330 , n11331 , n11332 , n11333 , n11336 , n11337 , n11338 , n11339 , n11342 , n11343 , n11344 , n11345 , n11348 , n11349 , n11350 , n11351 , n11354 , n11355 , n11356 , n11357 , n11360 , n11361 , n11362 , n11363 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11384 , n11385 , n11386 , n11387 , n11390 , n11391 , n11392 , n11393 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11422 , n11423 , n11424 , n11429 , n11430 , n11431 , n11432 , n11435 , n11436 , n11437 , n11438 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 ;
  assign n1205 = x57 & ~x59 ;
  assign n1206 = n1205 ^ x59 ;
  assign n1288 = ~x56 & ~x62 ;
  assign n1289 = ~x55 & n1288 ;
  assign n1290 = ~n1206 & n1289 ;
  assign n1349 = x216 & ~x221 ;
  assign n1350 = ~x215 & n1349 ;
  assign n1347 = ~x215 & x221 ;
  assign n1348 = n1347 ^ x215 ;
  assign n1351 = n1350 ^ n1348 ;
  assign n1352 = ~x216 & x833 ;
  assign n1353 = ~x215 & ~x929 ;
  assign n1354 = n1352 & n1353 ;
  assign n1355 = n1354 ^ x215 ;
  assign n1363 = ~x221 & ~n1355 ;
  assign n1364 = x265 & n1363 ;
  assign n1365 = n1364 ^ x265 ;
  assign n1357 = n1354 ^ x265 ;
  assign n1366 = n1365 ^ n1357 ;
  assign n1367 = ~x332 & ~n1366 ;
  assign n1373 = n1347 & n1352 ;
  assign n1374 = n1373 ^ n1348 ;
  assign n1377 = n1367 & n1374 ;
  assign n1378 = ~x1144 & n1377 ;
  assign n1379 = n1378 ^ x1144 ;
  assign n1368 = n1367 ^ x332 ;
  assign n1369 = n1368 ^ x1144 ;
  assign n1380 = n1379 ^ n1369 ;
  assign n1381 = n1351 & n1380 ;
  assign n1382 = ~n1290 & ~n1381 ;
  assign n1207 = ~x67 & ~x68 ;
  assign n1208 = ~x71 & ~x84 ;
  assign n1209 = n1207 & n1208 ;
  assign n1210 = ~x69 & ~x83 ;
  assign n1211 = ~x103 & n1210 ;
  assign n1212 = ~x66 & n1211 ;
  assign n1213 = x82 & ~x111 ;
  assign n1214 = n1213 ^ x111 ;
  assign n1215 = ~x36 & ~n1214 ;
  assign n1216 = ~x48 & ~x61 ;
  assign n1217 = ~x76 & ~x85 ;
  assign n1218 = ~x106 & n1217 ;
  assign n1219 = n1216 & n1218 ;
  assign n1221 = x104 & ~n1219 ;
  assign n1220 = n1219 ^ x104 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1223 = n1222 ^ x89 ;
  assign n1224 = ~x49 & ~n1221 ;
  assign n1225 = n1224 ^ x89 ;
  assign n1226 = ~n1223 & ~n1225 ;
  assign n1227 = n1226 ^ x89 ;
  assign n1228 = ~x45 & ~n1227 ;
  assign n1229 = ~x49 & ~x89 ;
  assign n1230 = n1222 & n1229 ;
  assign n1232 = ~n1228 & ~n1230 ;
  assign n1231 = n1230 ^ n1228 ;
  assign n1233 = n1232 ^ n1231 ;
  assign n1234 = n1215 & ~n1233 ;
  assign n1235 = n1212 & n1234 ;
  assign n1236 = ~x73 & n1235 ;
  assign n1237 = ~x81 & n1236 ;
  assign n1238 = ~x64 & ~x65 ;
  assign n1239 = ~x88 & ~x98 ;
  assign n1240 = ~x102 & ~x107 ;
  assign n1241 = n1239 & n1240 ;
  assign n1242 = ~x63 & n1241 ;
  assign n1243 = n1238 & n1242 ;
  assign n1244 = n1237 & n1243 ;
  assign n1245 = n1209 & n1244 ;
  assign n1246 = ~x53 & x60 ;
  assign n1247 = n1246 ^ x53 ;
  assign n1248 = ~x58 & ~n1247 ;
  assign n1250 = x97 & x108 ;
  assign n1249 = x108 ^ x97 ;
  assign n1251 = n1250 ^ n1249 ;
  assign n1252 = ~x94 & ~n1251 ;
  assign n1253 = ~x50 & ~x110 ;
  assign n1254 = ~x91 & ~x109 ;
  assign n1255 = ~x46 & ~x47 ;
  assign n1256 = n1254 & n1255 ;
  assign n1257 = ~x77 & ~x86 ;
  assign n1258 = n1256 & n1257 ;
  assign n1259 = n1253 & n1258 ;
  assign n1260 = n1252 & n1259 ;
  assign n1261 = n1248 & n1260 ;
  assign n1262 = n1245 & n1261 ;
  assign n1263 = ~x72 & ~x96 ;
  assign n1264 = ~x51 & ~x70 ;
  assign n1265 = n1263 & n1264 ;
  assign n1266 = x35 & ~x93 ;
  assign n1267 = n1266 ^ x93 ;
  assign n1268 = ~x90 & ~n1267 ;
  assign n1269 = n1265 & n1268 ;
  assign n1270 = n1262 & n1269 ;
  assign n1271 = ~x32 & ~x95 ;
  assign n1272 = ~x40 & n1271 ;
  assign n1273 = n1270 & n1272 ;
  assign n1291 = n1273 & n1290 ;
  assign n1277 = ~x38 & ~x54 ;
  assign n1292 = ~x74 & ~x75 ;
  assign n1293 = n1277 & n1292 ;
  assign n1294 = x92 ^ x87 ;
  assign n1295 = n1294 ^ x100 ;
  assign n1296 = n1295 ^ x39 ;
  assign n1297 = n1293 & n1296 ;
  assign n1298 = x92 ^ x39 ;
  assign n1299 = x100 ^ x92 ;
  assign n1300 = n1298 & n1299 ;
  assign n1301 = n1300 ^ x92 ;
  assign n1302 = n1297 & ~n1301 ;
  assign n1303 = n1291 & n1302 ;
  assign n1285 = x62 ^ x56 ;
  assign n1274 = ~x75 & x100 ;
  assign n1275 = n1274 ^ x75 ;
  assign n1276 = ~x87 & ~n1275 ;
  assign n1278 = ~x74 & ~x92 ;
  assign n1279 = n1277 & n1278 ;
  assign n1280 = n1276 & n1279 ;
  assign n1281 = x39 & n1280 ;
  assign n1282 = n1281 ^ n1280 ;
  assign n1283 = n1273 & n1282 ;
  assign n1284 = ~n1206 & n1283 ;
  assign n1286 = ~x55 & n1284 ;
  assign n1287 = n1285 & n1286 ;
  assign n1304 = n1303 ^ n1287 ;
  assign n1310 = ~x39 & ~x87 ;
  assign n1311 = ~x38 & n1310 ;
  assign n1312 = ~x92 & ~n1275 ;
  assign n1313 = n1311 & n1312 ;
  assign n1314 = ~x74 & n1313 ;
  assign n1315 = n1273 & n1314 ;
  assign n1316 = ~x57 & n1288 ;
  assign n1318 = ~x54 & ~x59 ;
  assign n1317 = x59 ^ x54 ;
  assign n1319 = n1318 ^ n1317 ;
  assign n1320 = n1316 & n1319 ;
  assign n1321 = n1318 ^ x55 ;
  assign n1322 = n1320 & ~n1321 ;
  assign n1323 = n1315 & n1322 ;
  assign n1305 = x38 & ~x39 ;
  assign n1306 = ~x54 & n1278 ;
  assign n1307 = n1276 & n1306 ;
  assign n1308 = n1291 & n1307 ;
  assign n1309 = n1305 & n1308 ;
  assign n1324 = n1323 ^ n1309 ;
  assign n1325 = n1283 & n1288 ;
  assign n1326 = n1205 & n1325 ;
  assign n1327 = ~x55 & n1326 ;
  assign n1328 = n1291 & n1311 ;
  assign n1329 = x74 ^ x54 ;
  assign n1330 = n1329 ^ x75 ;
  assign n1331 = n1330 ^ x92 ;
  assign n1332 = x75 ^ x74 ;
  assign n1333 = x92 ^ x74 ;
  assign n1334 = n1332 & n1333 ;
  assign n1335 = n1334 ^ x74 ;
  assign n1336 = n1331 & ~n1335 ;
  assign n1337 = n1328 & n1336 ;
  assign n1338 = ~x100 & n1337 ;
  assign n1339 = ~n1327 & ~n1338 ;
  assign n1340 = ~n1324 & n1339 ;
  assign n1341 = ~n1304 & n1340 ;
  assign n1344 = ~x105 & x228 ;
  assign n1345 = n1344 ^ x228 ;
  assign n1346 = x153 & ~n1345 ;
  assign n1383 = ~x137 & ~n1351 ;
  assign n1384 = ~n1344 & n1383 ;
  assign n1385 = n1384 ^ n1351 ;
  assign n1386 = n1346 & ~n1385 ;
  assign n1394 = ~n1206 & n1386 ;
  assign n1395 = ~x228 & n1394 ;
  assign n1396 = n1395 ^ x228 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1388 = n1387 ^ x228 ;
  assign n1397 = n1396 ^ n1388 ;
  assign n1398 = ~n1341 & ~n1397 ;
  assign n1399 = n1382 & ~n1398 ;
  assign n1342 = n1284 & ~n1341 ;
  assign n1404 = x95 & ~x479 ;
  assign n1405 = x234 & n1404 ;
  assign n1408 = ~n1342 & ~n1405 ;
  assign n1409 = n1345 & n1408 ;
  assign n1410 = n1409 ^ n1345 ;
  assign n1400 = n1345 ^ n1287 ;
  assign n1411 = n1410 ^ n1400 ;
  assign n1412 = ~n1351 & ~n1411 ;
  assign n1413 = n1399 & n1412 ;
  assign n1416 = n1413 ^ n1399 ;
  assign n1343 = ~x228 & n1342 ;
  assign n1414 = n1346 & n1413 ;
  assign n1415 = ~n1343 & n1414 ;
  assign n1417 = n1416 ^ n1415 ;
  assign n1527 = x224 ^ x222 ;
  assign n1530 = x833 & x929 ;
  assign n1531 = n1530 ^ x265 ;
  assign n1532 = ~x224 & n1531 ;
  assign n1533 = n1532 ^ x265 ;
  assign n1534 = n1527 & n1533 ;
  assign n1535 = n1534 ^ x222 ;
  assign n1536 = ~x223 & ~n1535 ;
  assign n1537 = ~x299 & n1290 ;
  assign n1538 = ~n1536 & n1537 ;
  assign n1545 = ~x224 & x833 ;
  assign n1546 = x222 & ~x223 ;
  assign n1547 = ~n1545 & n1546 ;
  assign n1548 = n1547 ^ x223 ;
  assign n1551 = n1538 & n1548 ;
  assign n1552 = x1144 & n1551 ;
  assign n1553 = n1552 ^ x1144 ;
  assign n1418 = ~n1282 & n1290 ;
  assign n1419 = ~x223 & ~x299 ;
  assign n1422 = x224 & n1419 ;
  assign n1420 = x222 & n1419 ;
  assign n1421 = ~x224 & n1420 ;
  assign n1423 = n1422 ^ n1421 ;
  assign n1424 = n1423 ^ n1419 ;
  assign n1425 = ~x137 & ~x332 ;
  assign n1426 = n1424 & n1425 ;
  assign n1427 = x299 & ~n1381 ;
  assign n1428 = ~x332 & ~n1385 ;
  assign n1436 = x153 & n1428 ;
  assign n1437 = n1344 & n1436 ;
  assign n1438 = n1437 ^ n1344 ;
  assign n1429 = n1428 ^ x332 ;
  assign n1430 = n1429 ^ n1344 ;
  assign n1439 = n1438 ^ n1430 ;
  assign n1440 = n1427 & ~n1439 ;
  assign n1441 = ~n1426 & ~n1440 ;
  assign n1442 = ~x39 & ~n1280 ;
  assign n1508 = ~x215 & x299 ;
  assign n1509 = n1349 ^ x221 ;
  assign n1510 = n1508 & n1509 ;
  assign n1511 = n1510 ^ n1508 ;
  assign n1444 = n1346 & n1511 ;
  assign n1445 = ~x332 & n1444 ;
  assign n1446 = n1511 ^ n1445 ;
  assign n1447 = n1446 ^ n1427 ;
  assign n1456 = n1307 & ~n1447 ;
  assign n1448 = ~x74 & ~n1275 ;
  assign n1449 = ~n1277 & n1448 ;
  assign n1450 = n1449 ^ n1448 ;
  assign n1451 = n1294 & n1450 ;
  assign n1457 = n1456 ^ n1451 ;
  assign n1458 = n1442 & n1457 ;
  assign n1459 = n1458 ^ n1280 ;
  assign n1460 = n1441 & n1459 ;
  assign n1461 = n1273 & n1460 ;
  assign n1462 = n1418 & ~n1461 ;
  assign n1463 = n1425 & n1427 ;
  assign n1464 = x137 & ~n1275 ;
  assign n1465 = x100 ^ x75 ;
  assign n1466 = n1306 & n1465 ;
  assign n1467 = ~x144 & ~x174 ;
  assign n1468 = ~x189 & n1467 ;
  assign n1469 = ~x198 & n1426 ;
  assign n1470 = ~x142 & n1469 ;
  assign n1471 = ~n1468 & n1470 ;
  assign n1472 = n1471 ^ n1469 ;
  assign n1473 = n1472 ^ n1426 ;
  assign n1474 = n1466 & ~n1473 ;
  assign n1475 = n1336 & ~n1474 ;
  assign n1476 = n1464 & n1475 ;
  assign n1477 = n1476 ^ n1474 ;
  assign n1478 = n1463 & n1477 ;
  assign n1482 = ~x152 & ~x161 ;
  assign n1483 = ~x166 & n1482 ;
  assign n1484 = ~x146 & ~n1483 ;
  assign n1489 = n1478 & ~n1484 ;
  assign n1490 = ~x210 & n1489 ;
  assign n1491 = n1490 ^ x210 ;
  assign n1479 = n1478 ^ n1477 ;
  assign n1480 = n1479 ^ x210 ;
  assign n1492 = n1491 ^ n1480 ;
  assign n1493 = n1273 & n1492 ;
  assign n1494 = n1311 & n1493 ;
  assign n1495 = n1494 ^ n1447 ;
  assign n1496 = ~x228 & n1273 ;
  assign n1497 = n1302 & n1496 ;
  assign n1498 = ~x39 & x252 ;
  assign n1499 = ~n1451 & n1498 ;
  assign n1500 = ~n1484 & n1499 ;
  assign n1501 = n1497 & n1500 ;
  assign n1502 = n1501 ^ n1497 ;
  assign n1503 = ~n1351 & n1502 ;
  assign n1504 = ~n1494 & n1503 ;
  assign n1505 = n1504 ^ n1494 ;
  assign n1512 = n1345 & n1511 ;
  assign n1513 = n1512 ^ n1424 ;
  assign n1518 = ~n1405 & n1513 ;
  assign n1519 = ~x332 & n1518 ;
  assign n1520 = n1519 ^ x332 ;
  assign n1506 = n1504 ^ x332 ;
  assign n1521 = n1520 ^ n1506 ;
  assign n1522 = ~n1505 & n1521 ;
  assign n1523 = n1522 ^ n1503 ;
  assign n1524 = ~n1495 & ~n1523 ;
  assign n1525 = n1524 ^ n1494 ;
  assign n1526 = n1462 & ~n1525 ;
  assign n1540 = n1538 ^ n1526 ;
  assign n1541 = n1540 ^ x1144 ;
  assign n1554 = n1553 ^ n1541 ;
  assign n1555 = ~n1417 & ~n1554 ;
  assign n1556 = n1418 ^ n1290 ;
  assign n1765 = ~x40 & x95 ;
  assign n1763 = x40 ^ x32 ;
  assign n1557 = ~x90 & n1262 ;
  assign n1558 = x93 ^ x35 ;
  assign n1559 = n1557 & n1558 ;
  assign n1560 = x110 ^ x90 ;
  assign n1561 = x90 ^ x58 ;
  assign n1562 = n1560 & ~n1561 ;
  assign n1563 = n1562 ^ x110 ;
  assign n1564 = x91 ^ x47 ;
  assign n1565 = ~x58 & ~x90 ;
  assign n1566 = n1565 ^ x91 ;
  assign n1567 = n1564 & ~n1566 ;
  assign n1568 = n1567 ^ x91 ;
  assign n1569 = ~n1267 & ~n1568 ;
  assign n1570 = n1567 ^ n1563 ;
  assign n1571 = n1570 ^ n1569 ;
  assign n1572 = n1567 ^ n1562 ;
  assign n1573 = n1572 ^ n1569 ;
  assign n1574 = n1562 ^ x47 ;
  assign n1575 = n1574 ^ n1563 ;
  assign n1576 = ~n1573 & n1575 ;
  assign n1577 = n1571 & n1576 ;
  assign n1578 = n1577 ^ n1562 ;
  assign n1579 = n1578 ^ n1563 ;
  assign n1580 = n1569 & ~n1579 ;
  assign n1581 = ~n1563 & n1580 ;
  assign n1582 = ~x50 & ~n1247 ;
  assign n1583 = ~x77 & n1582 ;
  assign n1584 = ~n1251 & n1583 ;
  assign n1586 = x86 & x94 ;
  assign n1585 = x94 ^ x86 ;
  assign n1587 = n1586 ^ n1585 ;
  assign n1588 = n1584 & ~n1587 ;
  assign n1589 = n1245 & n1588 ;
  assign n1590 = x46 & ~x109 ;
  assign n1591 = n1590 ^ x109 ;
  assign n1592 = x53 ^ x50 ;
  assign n1593 = n1592 ^ n1246 ;
  assign n1594 = n1247 ^ x60 ;
  assign n1595 = n1594 ^ n1246 ;
  assign n1596 = n1595 ^ n1247 ;
  assign n1599 = ~x77 & ~n1596 ;
  assign n1600 = n1599 ^ n1247 ;
  assign n1601 = n1593 & n1600 ;
  assign n1602 = n1601 ^ x50 ;
  assign n1603 = ~n1591 & ~n1602 ;
  assign n1604 = n1589 & n1603 ;
  assign n1605 = ~x47 & ~x110 ;
  assign n1606 = n1565 & n1605 ;
  assign n1607 = ~x91 & ~x93 ;
  assign n1608 = n1606 & n1607 ;
  assign n1609 = ~n1604 & ~n1608 ;
  assign n1610 = n1581 & n1609 ;
  assign n1611 = n1610 ^ n1581 ;
  assign n1739 = ~x46 & ~n1254 ;
  assign n1612 = n1583 ^ n1251 ;
  assign n1613 = ~n1250 & ~n1587 ;
  assign n1614 = n1613 ^ n1251 ;
  assign n1615 = ~n1612 & ~n1614 ;
  assign n1616 = n1615 ^ n1251 ;
  assign n1617 = n1245 & ~n1616 ;
  assign n1618 = n1588 & ~n1617 ;
  assign n1621 = n1209 & n1236 ;
  assign n1637 = ~x102 & n1209 ;
  assign n1638 = ~x81 & n1239 ;
  assign n1639 = n1637 & n1638 ;
  assign n1641 = n1639 ^ x63 ;
  assign n1624 = x98 ^ x88 ;
  assign n1625 = n1624 ^ x102 ;
  assign n1626 = n1625 ^ x107 ;
  assign n1627 = x102 ^ x98 ;
  assign n1629 = ~n1624 & n1627 ;
  assign n1630 = n1629 ^ x102 ;
  assign n1631 = n1626 & ~n1630 ;
  assign n1632 = n1631 ^ n1241 ;
  assign n1633 = ~x81 & n1632 ;
  assign n1634 = n1633 ^ n1241 ;
  assign n1642 = n1641 ^ n1634 ;
  assign n1622 = x65 ^ x64 ;
  assign n1623 = x65 ^ x63 ;
  assign n1635 = n1634 ^ n1623 ;
  assign n1636 = ~n1622 & n1635 ;
  assign n1640 = n1639 ^ n1636 ;
  assign n1643 = n1642 ^ n1640 ;
  assign n1644 = n1621 & ~n1643 ;
  assign n1649 = n1634 & n1640 ;
  assign n1650 = n1649 ^ n1639 ;
  assign n1651 = n1644 & n1650 ;
  assign n1654 = x68 ^ x66 ;
  assign n1655 = n1654 ^ x73 ;
  assign n1656 = n1655 ^ x84 ;
  assign n1657 = x73 ^ x68 ;
  assign n1658 = x84 ^ x73 ;
  assign n1659 = n1657 & ~n1658 ;
  assign n1660 = n1659 ^ x68 ;
  assign n1661 = ~x66 & ~n1660 ;
  assign n1662 = ~n1656 & n1661 ;
  assign n1663 = x106 ^ x85 ;
  assign n1664 = x85 ^ x76 ;
  assign n1665 = n1663 & n1664 ;
  assign n1666 = n1665 ^ x85 ;
  assign n1667 = n1216 & ~n1666 ;
  assign n1668 = n1667 ^ x48 ;
  assign n1669 = n1668 ^ x61 ;
  assign n1670 = n1669 ^ n1667 ;
  assign n1673 = n1218 & n1670 ;
  assign n1674 = n1673 ^ n1667 ;
  assign n1675 = n1662 & n1674 ;
  assign n1676 = ~n1232 & n1675 ;
  assign n1677 = ~n1233 & ~n1660 ;
  assign n1678 = n1656 & n1677 ;
  assign n1679 = ~n1676 & ~n1678 ;
  assign n1680 = ~n1233 & n1662 ;
  assign n1681 = n1211 & n1680 ;
  assign n1682 = x82 ^ x36 ;
  assign n1684 = x82 ^ x67 ;
  assign n1683 = x111 ^ x82 ;
  assign n1685 = n1684 ^ n1683 ;
  assign n1686 = n1685 ^ x82 ;
  assign n1687 = ~n1682 & n1686 ;
  assign n1688 = n1687 ^ n1685 ;
  assign n1689 = n1681 & ~n1688 ;
  assign n1698 = x111 & ~n1687 ;
  assign n1692 = n1689 ^ n1211 ;
  assign n1690 = ~x36 & ~x67 ;
  assign n1691 = ~n1214 & n1690 ;
  assign n1693 = n1692 ^ n1691 ;
  assign n1699 = n1698 ^ n1693 ;
  assign n1700 = n1689 & n1699 ;
  assign n1701 = n1700 ^ n1693 ;
  assign n1702 = n1701 ^ n1211 ;
  assign n1703 = n1701 ^ n1689 ;
  assign n1704 = ~n1700 & ~n1703 ;
  assign n1705 = ~n1702 & n1704 ;
  assign n1706 = n1705 ^ n1701 ;
  assign n1707 = ~n1679 & ~n1706 ;
  assign n1716 = ~x71 & ~x81 ;
  assign n1717 = n1243 & n1716 ;
  assign n1709 = n1680 & n1691 ;
  assign n1710 = n1709 ^ n1707 ;
  assign n1711 = x103 ^ x83 ;
  assign n1712 = x83 ^ x69 ;
  assign n1713 = n1711 & n1712 ;
  assign n1714 = n1713 ^ x83 ;
  assign n1715 = n1710 & ~n1714 ;
  assign n1720 = n1717 ^ n1715 ;
  assign n1721 = ~n1707 & ~n1720 ;
  assign n1708 = n1707 ^ n1244 ;
  assign n1722 = n1721 ^ n1708 ;
  assign n1723 = n1721 ^ n1709 ;
  assign n1718 = n1717 ^ n1707 ;
  assign n1724 = n1721 ^ n1718 ;
  assign n1725 = n1724 ^ n1707 ;
  assign n1726 = n1723 & ~n1725 ;
  assign n1727 = ~n1722 & n1726 ;
  assign n1728 = n1727 ^ n1724 ;
  assign n1731 = ~n1651 & n1728 ;
  assign n1732 = n1618 & n1731 ;
  assign n1733 = n1732 ^ n1618 ;
  assign n1734 = n1733 ^ n1617 ;
  assign n1735 = n1603 & n1734 ;
  assign n1736 = ~n1586 & n1735 ;
  assign n1740 = n1739 ^ n1736 ;
  assign n1741 = n1589 & n1740 ;
  assign n1742 = n1741 ^ n1736 ;
  assign n1743 = n1606 & n1742 ;
  assign n1744 = n1743 ^ n1606 ;
  assign n1745 = n1611 & ~n1744 ;
  assign n1746 = n1265 & n1272 ;
  assign n1747 = x96 ^ x51 ;
  assign n1748 = x72 ^ x70 ;
  assign n1749 = n1748 ^ x96 ;
  assign n1750 = ~n1747 & n1749 ;
  assign n1751 = n1750 ^ n1748 ;
  assign n1752 = n1262 & n1268 ;
  assign n1753 = n1272 & n1752 ;
  assign n1754 = ~n1751 & n1753 ;
  assign n1755 = x72 & ~n1750 ;
  assign n1756 = n1754 & n1755 ;
  assign n1757 = n1756 ^ n1754 ;
  assign n1758 = n1746 & ~n1757 ;
  assign n1759 = ~n1745 & n1758 ;
  assign n1760 = ~n1559 & n1759 ;
  assign n1761 = n1760 ^ n1758 ;
  assign n1762 = n1761 ^ n1757 ;
  assign n1764 = n1763 ^ n1762 ;
  assign n1766 = n1765 ^ n1764 ;
  assign n1767 = n1766 ^ n1762 ;
  assign n1768 = n1766 ^ x95 ;
  assign n1769 = n1768 ^ n1765 ;
  assign n1770 = n1769 ^ n1766 ;
  assign n1771 = n1767 & n1770 ;
  assign n1772 = n1771 ^ n1766 ;
  assign n1773 = n1270 & n1772 ;
  assign n1774 = n1773 ^ n1762 ;
  assign n1775 = ~x228 & n1774 ;
  assign n1776 = n1775 ^ n1345 ;
  assign n1777 = n1511 & n1776 ;
  assign n1778 = n1777 ^ n1424 ;
  assign n1782 = x210 ^ x198 ;
  assign n1783 = x299 & n1782 ;
  assign n1784 = n1783 ^ x198 ;
  assign n1785 = ~x841 & n1784 ;
  assign n1786 = n1785 ^ x841 ;
  assign n1787 = x225 & n1786 ;
  assign n1779 = ~x40 & n1270 ;
  assign n2734 = ~x70 & ~x95 ;
  assign n2735 = ~n1247 & n2734 ;
  assign n2736 = x32 & n2735 ;
  assign n2737 = n1779 & n2736 ;
  assign n1788 = n1787 & n2737 ;
  assign n1789 = n1778 & ~n1788 ;
  assign n1790 = ~n1746 & ~n1774 ;
  assign n1791 = n1483 ^ n1468 ;
  assign n1792 = x299 & n1791 ;
  assign n1793 = n1792 ^ n1468 ;
  assign n1794 = x146 ^ x142 ;
  assign n1795 = x299 & n1794 ;
  assign n1796 = n1795 ^ x142 ;
  assign n1797 = ~n1793 & ~n1796 ;
  assign n1798 = ~n1784 & ~n1797 ;
  assign n1799 = ~x40 & ~x51 ;
  assign n1800 = n1263 & n1799 ;
  assign n1801 = n1800 ^ x225 ;
  assign n1802 = ~x35 & n1801 ;
  assign n1803 = n1802 ^ x225 ;
  assign n1805 = n1557 ^ x93 ;
  assign n1806 = n1803 & n1805 ;
  assign n1807 = n1806 ^ x35 ;
  assign n1808 = n1557 & ~n1807 ;
  assign n1809 = ~x95 & ~n1808 ;
  assign n1810 = n1604 & n1605 ;
  assign n1811 = n1565 & n1589 ;
  assign n1812 = ~n1810 & n1811 ;
  assign n1816 = ~x109 & ~x110 ;
  assign n1821 = n1812 & ~n1816 ;
  assign n1822 = ~n1255 & n1821 ;
  assign n1823 = n1822 ^ n1255 ;
  assign n1813 = n1812 ^ n1565 ;
  assign n1814 = n1813 ^ n1255 ;
  assign n1824 = n1823 ^ n1814 ;
  assign n1825 = n1611 & ~n1824 ;
  assign n1826 = n1809 & ~n1825 ;
  assign n1827 = ~n1745 & n1826 ;
  assign n1828 = ~x97 & ~x137 ;
  assign n1836 = ~x35 & n1828 ;
  assign n1837 = ~n1247 & n1836 ;
  assign n1838 = n1837 ^ n1247 ;
  assign n1829 = n1828 ^ x137 ;
  assign n1830 = n1829 ^ n1247 ;
  assign n1839 = n1838 ^ n1830 ;
  assign n1840 = ~n1827 & ~n1839 ;
  assign n1844 = x950 & x1092 ;
  assign n1845 = x829 & n1844 ;
  assign n1846 = x1091 & x1093 ;
  assign n1848 = ~x833 & x957 ;
  assign n1849 = n1846 & n1848 ;
  assign n1847 = n1846 ^ x1093 ;
  assign n1850 = n1849 ^ n1847 ;
  assign n1851 = n1845 & ~n1850 ;
  assign n1852 = ~x841 & n1851 ;
  assign n1853 = x96 & n1757 ;
  assign n1869 = n1852 & n1853 ;
  assign n1854 = ~x35 & n1608 ;
  assign n1855 = n1746 & n1854 ;
  assign n1856 = x97 & n1608 ;
  assign n1857 = n1735 & n1856 ;
  assign n1858 = n1855 & n1857 ;
  assign n1860 = n1858 ^ n1853 ;
  assign n1861 = ~x46 & ~x94 ;
  assign n1862 = x97 ^ x36 ;
  assign n1863 = ~x1093 & n1845 ;
  assign n1864 = n1863 ^ n1851 ;
  assign n1865 = n1862 & n1864 ;
  assign n1866 = n1861 & n1865 ;
  assign n1867 = n1860 & ~n1866 ;
  assign n1870 = n1869 ^ n1867 ;
  assign n1871 = n1870 ^ n1860 ;
  assign n1876 = n1840 & n1871 ;
  assign n1877 = n1798 & n1876 ;
  assign n1878 = n1877 ^ n1798 ;
  assign n1841 = n1840 ^ n1827 ;
  assign n1842 = n1841 ^ n1798 ;
  assign n1879 = n1878 ^ n1842 ;
  assign n1880 = ~n1790 & ~n1879 ;
  assign n1881 = n1880 ^ x234 ;
  assign n1882 = ~n1404 & ~n1853 ;
  assign n1885 = n1881 & n1882 ;
  assign n1886 = n1885 ^ x234 ;
  assign n1887 = n1789 & ~n1886 ;
  assign n1888 = n1556 & n1887 ;
  assign n1889 = n1888 ^ n1556 ;
  assign n1892 = ~n1351 & n1776 ;
  assign n1897 = n1447 & ~n1892 ;
  assign n1898 = n1889 & n1897 ;
  assign n1899 = n1898 ^ n1889 ;
  assign n1900 = n1899 ^ n1556 ;
  assign n1901 = n1555 & ~n1900 ;
  assign n1902 = ~x332 & ~n1901 ;
  assign n1904 = ~n1345 & ~n1351 ;
  assign n1910 = n1904 ^ n1351 ;
  assign n1911 = ~n1404 & ~n1910 ;
  assign n1912 = n1911 ^ n1910 ;
  assign n1913 = x239 & ~n1912 ;
  assign n1909 = x939 & n1373 ;
  assign n1914 = n1913 ^ n1909 ;
  assign n1906 = x1146 & n1374 ;
  assign n1905 = ~x154 & n1904 ;
  assign n1907 = n1906 ^ n1905 ;
  assign n1903 = x276 & n1350 ;
  assign n1908 = n1907 ^ n1903 ;
  assign n1915 = n1914 ^ n1908 ;
  assign n1916 = ~n1351 & ~n1537 ;
  assign n1917 = n1290 & n1502 ;
  assign n1918 = n1916 & ~n1917 ;
  assign n1919 = n1556 & n1774 ;
  assign n1920 = ~n1342 & ~n1919 ;
  assign n1926 = ~x228 & ~n1920 ;
  assign n1921 = n1916 ^ n1537 ;
  assign n1927 = n1926 ^ n1921 ;
  assign n1928 = n1918 & n1927 ;
  assign n1929 = n1928 ^ n1921 ;
  assign n1930 = n1915 & ~n1929 ;
  assign n1935 = n1421 ^ n1420 ;
  assign n1936 = n1935 ^ n1422 ;
  assign n1937 = x276 & n1936 ;
  assign n1933 = ~x299 & n1548 ;
  assign n1934 = x1146 & n1933 ;
  assign n1938 = n1937 ^ n1934 ;
  assign n1931 = n1420 & n1545 ;
  assign n1932 = x939 & n1931 ;
  assign n1939 = n1938 ^ n1932 ;
  assign n1940 = n1290 & ~n1939 ;
  assign n1944 = n1775 & ~n1882 ;
  assign n1945 = n1282 & ~n1351 ;
  assign n1946 = x299 & n1945 ;
  assign n1947 = n1282 & ~n1404 ;
  assign n1948 = n1853 & n1947 ;
  assign n1949 = n1948 ^ n1404 ;
  assign n1950 = n1513 & n1949 ;
  assign n1951 = n1946 & ~n1950 ;
  assign n1952 = n1944 & n1951 ;
  assign n1953 = n1952 ^ n1950 ;
  assign n1958 = n1940 & n1953 ;
  assign n1959 = x239 & n1958 ;
  assign n1960 = n1959 ^ x239 ;
  assign n1941 = n1940 ^ n1290 ;
  assign n1942 = n1941 ^ x239 ;
  assign n1961 = n1960 ^ n1942 ;
  assign n1962 = ~n1930 & ~n1961 ;
  assign n1969 = x927 & n1373 ;
  assign n1968 = x235 & ~n1912 ;
  assign n1970 = n1969 ^ n1968 ;
  assign n1966 = ~x274 & n1350 ;
  assign n1964 = x1145 & n1374 ;
  assign n1963 = ~x151 & n1904 ;
  assign n1965 = n1964 ^ n1963 ;
  assign n1967 = n1966 ^ n1965 ;
  assign n1971 = n1970 ^ n1967 ;
  assign n1972 = ~n1929 & n1971 ;
  assign n1975 = ~x274 & n1936 ;
  assign n1974 = x1145 & n1933 ;
  assign n1976 = n1975 ^ n1974 ;
  assign n1973 = x927 & n1931 ;
  assign n1977 = n1976 ^ n1973 ;
  assign n1978 = n1290 & ~n1977 ;
  assign n1986 = x235 & n1978 ;
  assign n1987 = n1953 & n1986 ;
  assign n1988 = n1987 ^ n1953 ;
  assign n1979 = n1978 ^ n1290 ;
  assign n1980 = n1979 ^ n1953 ;
  assign n1989 = n1988 ^ n1980 ;
  assign n1990 = ~n1972 & ~n1989 ;
  assign n2045 = x284 & n1424 ;
  assign n2038 = ~x944 & n1290 ;
  assign n2039 = n1931 & n2038 ;
  assign n2040 = n2039 ^ n1936 ;
  assign n2041 = n2039 ^ n1290 ;
  assign n2042 = x264 & n2041 ;
  assign n2043 = n2040 & n2042 ;
  assign n2044 = n2043 ^ n2041 ;
  assign n2046 = ~n1949 & n2044 ;
  assign n2047 = n2045 & n2046 ;
  assign n2048 = n2047 ^ n2044 ;
  assign n2049 = ~x1143 & n1933 ;
  assign n2050 = n2048 & n2049 ;
  assign n2055 = n2050 ^ x238 ;
  assign n2021 = x284 & n1882 ;
  assign n2022 = n2021 ^ x146 ;
  assign n2023 = n1776 & ~n2022 ;
  assign n2024 = n2023 ^ x146 ;
  assign n2025 = n1945 & ~n2024 ;
  assign n2026 = n2025 ^ n1945 ;
  assign n1996 = x1143 & n1374 ;
  assign n1995 = x146 & n1904 ;
  assign n1997 = n1996 ^ n1995 ;
  assign n1994 = ~x284 & n1911 ;
  assign n1998 = n1997 ^ n1994 ;
  assign n1992 = x944 & n1373 ;
  assign n1991 = ~x264 & n1350 ;
  assign n1993 = n1992 ^ n1991 ;
  assign n1999 = n1998 ^ n1993 ;
  assign n2027 = x299 & ~n1503 ;
  assign n2028 = n1999 & n2027 ;
  assign n2000 = ~n1344 & ~n1351 ;
  assign n2001 = x284 & ~n1404 ;
  assign n2002 = n2000 & n2001 ;
  assign n2003 = n2002 ^ n2000 ;
  assign n2029 = n2028 ^ n2003 ;
  assign n2030 = n1502 ^ n1345 ;
  assign n2031 = n2028 ^ x299 ;
  assign n2032 = ~n1946 & n2031 ;
  assign n2033 = n2030 & n2032 ;
  assign n2034 = n2029 & n2033 ;
  assign n2035 = n2034 ^ n2032 ;
  assign n2036 = n2035 ^ n1946 ;
  assign n2037 = ~n2026 & n2036 ;
  assign n2051 = n2050 ^ n2048 ;
  assign n2052 = ~n2037 & n2051 ;
  assign n2056 = n1953 & n2052 ;
  assign n2057 = ~n2055 & n2056 ;
  assign n2004 = n2003 ^ n1999 ;
  assign n2012 = x238 & ~n1999 ;
  assign n2013 = x228 & n2012 ;
  assign n2014 = n2013 ^ x228 ;
  assign n2005 = n1343 & ~n1351 ;
  assign n2006 = n2005 ^ x228 ;
  assign n2015 = n2014 ^ n2006 ;
  assign n2016 = n2004 & ~n2015 ;
  assign n2017 = n2016 ^ n2003 ;
  assign n2018 = ~n1290 & n2017 ;
  assign n2054 = n2052 ^ n2018 ;
  assign n2058 = n2057 ^ n2054 ;
  assign n2068 = x216 & ~x277 ;
  assign n2061 = x1142 ^ x932 ;
  assign n2062 = ~n1352 & n2061 ;
  assign n2063 = n2062 ^ x932 ;
  assign n2069 = n2068 ^ n2063 ;
  assign n2070 = ~x221 & n2069 ;
  assign n2071 = n2070 ^ n2063 ;
  assign n2072 = n1508 & ~n2071 ;
  assign n2059 = ~x249 & ~n1882 ;
  assign n2060 = n1424 & n2059 ;
  assign n2073 = n2072 ^ n2060 ;
  assign n2074 = n1556 & n2073 ;
  assign n2075 = ~x249 & n1404 ;
  assign n2076 = ~n1910 & n2075 ;
  assign n2110 = ~x172 & ~n1343 ;
  assign n2111 = n2110 ^ n1404 ;
  assign n2112 = ~n1345 & n2111 ;
  assign n2113 = n2112 ^ n1404 ;
  assign n2114 = ~x262 & ~n2113 ;
  assign n2118 = n1345 ^ n1343 ;
  assign n2123 = n2114 & ~n2118 ;
  assign n2124 = ~n1917 & n2123 ;
  assign n2125 = n2124 ^ n1917 ;
  assign n2115 = n2114 ^ n2113 ;
  assign n2116 = n2115 ^ n1917 ;
  assign n2126 = n2125 ^ n2116 ;
  assign n2127 = ~n1351 & n2126 ;
  assign n2128 = n2071 ^ x1142 ;
  assign n2131 = ~x215 & n2128 ;
  assign n2132 = n2131 ^ x1142 ;
  assign n2133 = ~n2127 & ~n2132 ;
  assign n2134 = n2133 ^ n1503 ;
  assign n2135 = n2134 ^ n1290 ;
  assign n2136 = n1503 ^ x299 ;
  assign n2137 = n2136 ^ n1290 ;
  assign n2138 = x299 ^ x262 ;
  assign n2139 = n2138 ^ n2133 ;
  assign n2140 = n2137 & ~n2139 ;
  assign n2141 = ~n2135 & n2140 ;
  assign n2142 = n2141 ^ x299 ;
  assign n2143 = n2142 ^ n2133 ;
  assign n2144 = n1290 & ~n2143 ;
  assign n2145 = ~n2133 & n2144 ;
  assign n2146 = n2145 ^ n2133 ;
  assign n2151 = n2076 & ~n2146 ;
  assign n2087 = n1424 & ~n2075 ;
  assign n2101 = x262 & n2087 ;
  assign n2102 = ~n1949 & n2101 ;
  assign n2103 = n2102 ^ n1949 ;
  assign n2090 = ~x277 & n1936 ;
  assign n2089 = x1142 & n1933 ;
  assign n2091 = n2090 ^ n2089 ;
  assign n2088 = x932 & n1931 ;
  assign n2092 = n2091 ^ n2088 ;
  assign n2094 = n2092 ^ n2087 ;
  assign n2095 = n2094 ^ n1949 ;
  assign n2104 = n2103 ^ n2095 ;
  assign n2105 = n1290 & n2104 ;
  assign n2147 = ~n2105 & n2146 ;
  assign n2080 = x262 ^ x172 ;
  assign n2077 = x249 ^ x172 ;
  assign n2081 = n2080 ^ n2077 ;
  assign n2082 = n1882 & ~n2081 ;
  assign n2083 = n2082 ^ n2077 ;
  assign n2084 = n1776 & ~n2083 ;
  assign n2085 = n2084 ^ x172 ;
  assign n2086 = n1511 & ~n2085 ;
  assign n2148 = n2147 ^ n2086 ;
  assign n2152 = n2151 ^ n2148 ;
  assign n2153 = ~n2074 & ~n2152 ;
  assign n2154 = n2153 ^ n2086 ;
  assign n2155 = x241 & n1953 ;
  assign n2181 = x270 & n1936 ;
  assign n2180 = ~x1141 & n1933 ;
  assign n2182 = n2181 ^ n2180 ;
  assign n2179 = ~x935 & n1931 ;
  assign n2183 = n2182 ^ n2179 ;
  assign n2165 = x861 & ~n1404 ;
  assign n2185 = n2165 ^ x861 ;
  assign n2166 = n2165 ^ x171 ;
  assign n2169 = n1345 & ~n2166 ;
  assign n2170 = n2169 ^ x171 ;
  assign n2171 = ~n1351 & n2170 ;
  assign n2161 = ~x1141 & n1374 ;
  assign n2160 = x270 & n1350 ;
  assign n2162 = n2161 ^ n2160 ;
  assign n2159 = ~x935 & n1373 ;
  assign n2163 = n2162 ^ n2159 ;
  assign n2172 = n2171 ^ n2163 ;
  assign n2184 = n2172 ^ n2165 ;
  assign n2186 = n2185 ^ n2184 ;
  assign n2189 = ~n1503 & ~n2186 ;
  assign n2190 = n2189 ^ n2185 ;
  assign n2191 = x299 & n2190 ;
  assign n2192 = n2191 ^ n2165 ;
  assign n2193 = ~n1282 & n2192 ;
  assign n2194 = x299 & n1282 ;
  assign n2195 = ~n1892 & n2194 ;
  assign n2196 = n2172 & n2195 ;
  assign n2197 = n2196 ^ n2194 ;
  assign n2198 = n2197 ^ x299 ;
  assign n2199 = n1778 & ~n2198 ;
  assign n2206 = ~n1853 & n2165 ;
  assign n2207 = n2199 & n2206 ;
  assign n2208 = n2207 ^ n2199 ;
  assign n2209 = n2208 ^ n2198 ;
  assign n2210 = ~n2193 & n2209 ;
  assign n2211 = ~n2183 & ~n2210 ;
  assign n2212 = n1290 & ~n2211 ;
  assign n2215 = n2155 & n2212 ;
  assign n2156 = x241 & ~n1290 ;
  assign n2157 = ~n1912 & n2156 ;
  assign n2158 = n2157 ^ n1290 ;
  assign n2176 = ~n2005 & ~n2186 ;
  assign n2177 = n2176 ^ x861 ;
  assign n2178 = ~n2158 & ~n2177 ;
  assign n2213 = n2212 ^ n2178 ;
  assign n2216 = n2215 ^ n2213 ;
  assign n2217 = n2005 ^ n1911 ;
  assign n2222 = ~x1140 & n1374 ;
  assign n2221 = x282 & n1350 ;
  assign n2223 = n2222 ^ n2221 ;
  assign n2220 = ~x921 & n1373 ;
  assign n2224 = n2223 ^ n2220 ;
  assign n2219 = n1351 ^ x869 ;
  assign n2225 = n2224 ^ n2219 ;
  assign n2218 = ~x170 & n1904 ;
  assign n2226 = n2225 ^ n2218 ;
  assign n2227 = ~n2217 & n2226 ;
  assign n2228 = n2227 ^ x869 ;
  assign n2259 = x248 & ~n2228 ;
  assign n2260 = ~n1912 & n2259 ;
  assign n2261 = n2260 ^ n1912 ;
  assign n2229 = x299 & ~n2224 ;
  assign n2230 = x869 ^ x170 ;
  assign n2231 = n1282 & n1775 ;
  assign n2233 = n2231 ^ n2030 ;
  assign n2236 = ~n2230 & ~n2233 ;
  assign n2237 = n2236 ^ x869 ;
  assign n2238 = ~n1351 & ~n2237 ;
  assign n2239 = n2229 & ~n2238 ;
  assign n2245 = ~x282 & n1936 ;
  assign n2244 = x921 & n1931 ;
  assign n2246 = n2245 ^ n2244 ;
  assign n2242 = x1140 & n1933 ;
  assign n2240 = ~n1404 & n1424 ;
  assign n2241 = x869 & n2240 ;
  assign n2243 = n2242 ^ n2241 ;
  assign n2247 = n2246 ^ n2243 ;
  assign n2248 = ~n2239 & ~n2247 ;
  assign n2249 = n2248 ^ x248 ;
  assign n2250 = ~n1953 & ~n2249 ;
  assign n2251 = n2250 ^ x248 ;
  assign n2252 = n2251 ^ n2228 ;
  assign n2253 = n2252 ^ n1912 ;
  assign n2262 = n2261 ^ n2253 ;
  assign n2263 = ~n1290 & n2262 ;
  assign n2264 = n2263 ^ n2251 ;
  assign n2286 = x281 & n1350 ;
  assign n2285 = ~x1139 & n1374 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2283 = ~x920 & n1373 ;
  assign n2282 = x148 & n1904 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2288 = n2287 ^ n2284 ;
  assign n2292 = n2288 ^ x862 ;
  assign n2293 = n2292 ^ x247 ;
  assign n2294 = ~n1404 & n2293 ;
  assign n2295 = n2294 ^ x247 ;
  assign n2296 = ~n1910 & ~n2295 ;
  assign n2297 = n2296 ^ n2292 ;
  assign n2326 = ~n2005 & ~n2297 ;
  assign n2327 = n2326 ^ x862 ;
  assign n2328 = ~n1290 & n2327 ;
  assign n2314 = x862 ^ x247 ;
  assign n2270 = n1882 & n2314 ;
  assign n2265 = x247 ^ x148 ;
  assign n2271 = n2270 ^ n2265 ;
  assign n2272 = n1776 & ~n2271 ;
  assign n2273 = n2272 ^ x148 ;
  assign n2274 = n1946 & n2273 ;
  assign n2317 = ~n1949 & n2314 ;
  assign n2318 = n2317 ^ x247 ;
  assign n2490 = n1290 & n1424 ;
  assign n2319 = ~n2318 & n2490 ;
  assign n2275 = ~x920 & n1290 ;
  assign n2276 = n1931 & n2275 ;
  assign n2277 = n2276 ^ n1936 ;
  assign n2278 = n2276 ^ n1290 ;
  assign n2279 = x281 & n2278 ;
  assign n2280 = n2277 & n2279 ;
  assign n2281 = n2280 ^ n2278 ;
  assign n2307 = ~x1139 & n1548 ;
  assign n2298 = n2297 ^ x862 ;
  assign n2301 = ~n1945 & n2298 ;
  assign n2302 = n2301 ^ x862 ;
  assign n2303 = ~n1503 & ~n2302 ;
  assign n2304 = n2303 ^ x862 ;
  assign n2308 = n2307 ^ n2304 ;
  assign n2309 = ~x299 & ~n2308 ;
  assign n2310 = n2309 ^ n2304 ;
  assign n2311 = n2281 & ~n2310 ;
  assign n2312 = n2311 ^ n2281 ;
  assign n2320 = n2319 ^ n2312 ;
  assign n2321 = ~n2274 & n2320 ;
  assign n2329 = n2328 ^ n2321 ;
  assign n2346 = x877 & ~n1404 ;
  assign n2347 = n2346 ^ x169 ;
  assign n2375 = n2118 & ~n2347 ;
  assign n2376 = n2375 ^ x169 ;
  assign n2377 = ~n1351 & n2376 ;
  assign n2332 = x269 & n1350 ;
  assign n2331 = ~x1138 & n1374 ;
  assign n2333 = n2332 ^ n2331 ;
  assign n2330 = ~x940 & n1373 ;
  assign n2334 = n2333 ^ n2330 ;
  assign n2378 = n2377 ^ n2334 ;
  assign n2379 = ~n1290 & n2378 ;
  assign n2381 = x246 & ~n1912 ;
  assign n2382 = n2379 & n2381 ;
  assign n2335 = x299 & ~n2334 ;
  assign n2352 = n2030 & ~n2347 ;
  assign n2339 = x877 ^ x169 ;
  assign n2336 = x246 ^ x169 ;
  assign n2340 = n2339 ^ n2336 ;
  assign n2341 = n1882 & n2340 ;
  assign n2342 = n2341 ^ n2336 ;
  assign n2343 = n1776 & ~n2342 ;
  assign n2353 = n2352 ^ n2343 ;
  assign n2354 = ~n1282 & n2353 ;
  assign n2344 = n2343 ^ x169 ;
  assign n2355 = n2354 ^ n2344 ;
  assign n2356 = ~n1351 & n2355 ;
  assign n2357 = n2335 & ~n2356 ;
  assign n2361 = x940 & n1931 ;
  assign n2360 = ~x269 & n1936 ;
  assign n2362 = n2361 ^ n2360 ;
  assign n2363 = n2362 ^ x246 ;
  assign n2359 = x877 & n1424 ;
  assign n2364 = n2363 ^ n2359 ;
  assign n2358 = x1138 & n1933 ;
  assign n2365 = n2364 ^ n2358 ;
  assign n2366 = ~n1950 & n2365 ;
  assign n2367 = n2366 ^ x246 ;
  assign n2368 = n1290 & ~n2367 ;
  assign n2369 = ~n2357 & n2368 ;
  assign n2380 = n2379 ^ n2369 ;
  assign n2383 = n2382 ^ n2380 ;
  assign n2384 = x240 & n1424 ;
  assign n2386 = ~n1282 & ~n1950 ;
  assign n2385 = n1950 ^ n1282 ;
  assign n2387 = n2386 ^ n2385 ;
  assign n2389 = x933 & n1373 ;
  assign n2388 = x1137 & n1374 ;
  assign n2390 = n2389 ^ n2388 ;
  assign n2391 = x299 & ~n2390 ;
  assign n2399 = ~x280 & n1350 ;
  assign n2392 = x878 & ~n1404 ;
  assign n2393 = n2392 ^ x168 ;
  assign n2396 = n1345 & ~n2393 ;
  assign n2397 = n2396 ^ x168 ;
  assign n2398 = ~n1351 & ~n2397 ;
  assign n2401 = n2399 ^ n2398 ;
  assign n2402 = n2401 ^ x878 ;
  assign n2405 = ~n1503 & n2402 ;
  assign n2406 = n2405 ^ x878 ;
  assign n2407 = n2391 & ~n2406 ;
  assign n2408 = n2387 & ~n2407 ;
  assign n2409 = ~n1946 & n2408 ;
  assign n2410 = n1511 & ~n2386 ;
  assign n2414 = x878 ^ x168 ;
  assign n2411 = x240 ^ x168 ;
  assign n2415 = n2414 ^ n2411 ;
  assign n2416 = n1882 & n2415 ;
  assign n2417 = n2416 ^ n2411 ;
  assign n2418 = n1776 & ~n2417 ;
  assign n2419 = n2418 ^ x168 ;
  assign n2420 = n2410 & ~n2419 ;
  assign n2421 = ~n2409 & ~n2420 ;
  assign n2426 = ~x933 & n1931 ;
  assign n2425 = n1424 & ~n2392 ;
  assign n2427 = n2426 ^ n2425 ;
  assign n2423 = x280 & n1936 ;
  assign n2422 = ~x1137 & n1933 ;
  assign n2424 = n2423 ^ n2422 ;
  assign n2428 = n2427 ^ n2424 ;
  assign n2429 = ~n2421 & ~n2428 ;
  assign n2438 = n1949 & ~n2429 ;
  assign n2439 = n2384 & n2438 ;
  assign n2431 = n2390 ^ x878 ;
  assign n2432 = n2431 ^ n2401 ;
  assign n2430 = x240 & ~n1912 ;
  assign n2433 = n2432 ^ n2430 ;
  assign n2434 = ~n2005 & n2433 ;
  assign n2435 = n2434 ^ x878 ;
  assign n2436 = n2435 ^ n2429 ;
  assign n2440 = n2439 ^ n2436 ;
  assign n2441 = n1290 & n2440 ;
  assign n2442 = n2441 ^ n2435 ;
  assign n2445 = x266 & n1350 ;
  assign n2444 = x1136 & n1374 ;
  assign n2446 = n2445 ^ n2444 ;
  assign n2443 = x928 & n1373 ;
  assign n2447 = n2446 ^ n2443 ;
  assign n2448 = ~n1537 & ~n2447 ;
  assign n2449 = ~x875 & ~n1404 ;
  assign n2450 = n2449 ^ x166 ;
  assign n2453 = n2118 & ~n2450 ;
  assign n2454 = n2453 ^ x166 ;
  assign n2455 = ~n1556 & ~n2454 ;
  assign n2456 = n2455 ^ n1776 ;
  assign n2492 = x875 ^ x245 ;
  assign n2460 = n1882 & n2492 ;
  assign n2458 = n1290 ^ x245 ;
  assign n2461 = n2460 ^ n2458 ;
  assign n2462 = n2461 ^ n1290 ;
  assign n2463 = n1404 ^ x166 ;
  assign n2464 = n2463 ^ n2449 ;
  assign n2465 = n2030 & ~n2464 ;
  assign n2466 = n2465 ^ x166 ;
  assign n2469 = n2461 ^ n1418 ;
  assign n2470 = n2466 & ~n2469 ;
  assign n2471 = ~n2462 & n2470 ;
  assign n2472 = n2471 ^ n2462 ;
  assign n2473 = n2472 ^ n1290 ;
  assign n2474 = ~n2455 & ~n2473 ;
  assign n2475 = n2474 ^ n1290 ;
  assign n2476 = n2456 & ~n2475 ;
  assign n2477 = n2476 ^ n1776 ;
  assign n2478 = ~n1776 & ~n2466 ;
  assign n2479 = n1290 & n2478 ;
  assign n2480 = n2479 ^ n1351 ;
  assign n2481 = ~n1351 & ~n2480 ;
  assign n2482 = ~n2477 & n2481 ;
  assign n2483 = n2448 & ~n2482 ;
  assign n2495 = ~n1949 & n2492 ;
  assign n2496 = n2495 ^ x245 ;
  assign n2497 = n2490 & ~n2496 ;
  assign n2486 = ~x266 & n1936 ;
  assign n2485 = ~x1136 & n1933 ;
  assign n2487 = n2486 ^ n2485 ;
  assign n2484 = ~x928 & n1931 ;
  assign n2488 = n2487 ^ n2484 ;
  assign n2489 = n1290 & n2488 ;
  assign n2498 = n2497 ^ n2489 ;
  assign n2499 = ~n2483 & ~n2498 ;
  assign n2501 = x244 ^ x161 ;
  assign n2500 = x879 ^ x161 ;
  assign n2502 = n2501 ^ n2500 ;
  assign n2505 = ~n1404 & n2502 ;
  assign n2506 = n2505 ^ n2501 ;
  assign n2507 = n2118 & n2506 ;
  assign n2508 = n2507 ^ x161 ;
  assign n2509 = ~n1351 & n2508 ;
  assign n2510 = ~n1290 & ~n2509 ;
  assign n2511 = x938 & n1290 ;
  assign n2512 = n1931 & n2511 ;
  assign n2513 = n2512 ^ n1936 ;
  assign n2514 = n2512 ^ n1290 ;
  assign n2515 = x879 & ~n1949 ;
  assign n2520 = n1511 & n2030 ;
  assign n2521 = n2520 ^ n1424 ;
  assign n2522 = n2515 & n2521 ;
  assign n2523 = n2514 & ~n2522 ;
  assign n2524 = x279 & n2523 ;
  assign n2525 = n2513 & n2524 ;
  assign n2526 = n2525 ^ n2523 ;
  assign n2527 = n2526 ^ x244 ;
  assign n2528 = x1135 & n1933 ;
  assign n2529 = n2526 & n2528 ;
  assign n2530 = n2529 ^ n2526 ;
  assign n2531 = n1953 & n2530 ;
  assign n2532 = ~n2527 & n2531 ;
  assign n2533 = n2532 ^ n2530 ;
  assign n2534 = ~n1351 & n2533 ;
  assign n2535 = n2515 ^ x161 ;
  assign n2538 = ~n2233 & n2535 ;
  assign n2539 = n2538 ^ n2515 ;
  assign n2540 = n2534 & n2539 ;
  assign n2541 = n2540 ^ n2533 ;
  assign n2542 = ~n2510 & ~n2541 ;
  assign n2545 = x279 & n1350 ;
  assign n2544 = x1135 & n1374 ;
  assign n2546 = n2545 ^ n2544 ;
  assign n2543 = x938 & n1373 ;
  assign n2547 = n2546 ^ n2543 ;
  assign n2548 = ~n2542 & ~n2547 ;
  assign n2549 = ~x299 & n2533 ;
  assign n2550 = ~n2548 & n2549 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2563 = x846 ^ x242 ;
  assign n2557 = ~n1404 & n2563 ;
  assign n2552 = x242 ^ x152 ;
  assign n2558 = n2557 ^ n2552 ;
  assign n2559 = n2118 & n2558 ;
  assign n2560 = n2559 ^ x152 ;
  assign n2561 = ~n1351 & ~n2560 ;
  assign n2562 = ~n1290 & ~n2561 ;
  assign n2564 = ~n1949 & n2563 ;
  assign n2565 = n2564 ^ x242 ;
  assign n2566 = n1424 & ~n2565 ;
  assign n2568 = ~x278 & n1936 ;
  assign n2567 = ~x930 & n1931 ;
  assign n2569 = n2568 ^ n2567 ;
  assign n2570 = n1290 & ~n2569 ;
  assign n2571 = n2566 & n2570 ;
  assign n2572 = n2571 ^ n2570 ;
  assign n2573 = ~n1351 & n2572 ;
  assign n2574 = n2565 ^ x152 ;
  assign n2577 = ~n2233 & n2574 ;
  assign n2578 = n2577 ^ n2565 ;
  assign n2579 = n2573 & ~n2578 ;
  assign n2580 = n2579 ^ n2572 ;
  assign n2581 = ~n2562 & ~n2580 ;
  assign n2583 = ~x930 & n1373 ;
  assign n2582 = ~x278 & n1350 ;
  assign n2584 = n2583 ^ n2582 ;
  assign n2585 = ~n2581 & ~n2584 ;
  assign n2595 = ~x299 & n2572 ;
  assign n2589 = n2585 ^ x1134 ;
  assign n2586 = n1933 ^ n1374 ;
  assign n2587 = n1537 & n2586 ;
  assign n2588 = n2587 ^ n1374 ;
  assign n2590 = n2589 ^ n2588 ;
  assign n2596 = n2595 ^ n2590 ;
  assign n2597 = ~n2585 & n2596 ;
  assign n2598 = n2597 ^ n2590 ;
  assign n2599 = n2598 ^ x1134 ;
  assign n2600 = n2598 ^ n2585 ;
  assign n2601 = ~n2597 & n2600 ;
  assign n2602 = n2599 & n2601 ;
  assign n2603 = n2602 ^ n2598 ;
  assign n2717 = x93 & x841 ;
  assign n2718 = n1559 & n1800 ;
  assign n2719 = ~n2717 & n2718 ;
  assign n2720 = n2719 ^ n1800 ;
  assign n2721 = n1245 & n1252 ;
  assign n2722 = n1611 & ~n2721 ;
  assign n2723 = n1736 & n2722 ;
  assign n2724 = n2723 ^ n2720 ;
  assign n2725 = n2720 & n2724 ;
  assign n2726 = ~n1825 & n2725 ;
  assign n2727 = ~n1790 & ~n2726 ;
  assign n2728 = ~n1779 & ~n2727 ;
  assign n2729 = ~n1273 & n1556 ;
  assign n2730 = ~n2728 & n2729 ;
  assign n2733 = x32 & n2730 ;
  assign n2738 = n1786 & n2737 ;
  assign n2739 = n2738 ^ n2736 ;
  assign n2740 = n2739 ^ n2735 ;
  assign n2741 = n2733 & ~n2740 ;
  assign n2604 = n1327 ^ n1287 ;
  assign n2605 = ~x250 & n1797 ;
  assign n2606 = x824 & n1844 ;
  assign n2607 = ~x1093 & n2606 ;
  assign n2608 = ~n1863 & ~n2607 ;
  assign n2609 = n2605 & ~n2608 ;
  assign n2610 = ~x41 & ~x101 ;
  assign n2611 = ~x99 & n2610 ;
  assign n2612 = ~x113 & n2611 ;
  assign n2613 = ~x115 & ~x116 ;
  assign n2614 = ~x42 & ~x43 ;
  assign n2615 = ~x44 & ~x114 ;
  assign n2616 = n2614 & n2615 ;
  assign n2617 = n2613 & n2616 ;
  assign n2618 = n2612 & n2617 ;
  assign n2619 = ~x52 & n2618 ;
  assign n2620 = x683 & ~n2619 ;
  assign n2628 = ~x129 & n2620 ;
  assign n2629 = x250 & n2628 ;
  assign n2630 = n2629 ^ x250 ;
  assign n2621 = n2620 ^ x252 ;
  assign n2622 = n2621 ^ x250 ;
  assign n2631 = n2630 ^ n2622 ;
  assign n2632 = n1797 & n2631 ;
  assign n2633 = n2632 ^ x252 ;
  assign n2634 = n2609 & n2633 ;
  assign n2635 = n2634 ^ n2633 ;
  assign n2636 = n2635 ^ n1311 ;
  assign n2641 = ~x87 & x100 ;
  assign n2642 = n2636 & n2641 ;
  assign n2643 = n2642 ^ n2636 ;
  assign n2644 = n2643 ^ n2635 ;
  assign n2645 = ~x74 & n2644 ;
  assign n2646 = x39 & ~n2645 ;
  assign n2649 = ~x979 & ~x984 ;
  assign n2650 = ~x287 & n2649 ;
  assign n2651 = ~x252 & ~x1001 ;
  assign n2652 = x835 & ~n2651 ;
  assign n2653 = n2650 & n2652 ;
  assign n2654 = n1864 & n2653 ;
  assign n2674 = x299 & n1347 ;
  assign n2675 = ~x216 & n2674 ;
  assign n2676 = n2675 ^ n2674 ;
  assign n2655 = ~x332 & ~x468 ;
  assign n2677 = ~x970 & ~x972 ;
  assign n2678 = ~x975 & ~x978 ;
  assign n2679 = n2677 & n2678 ;
  assign n2680 = ~x907 & ~x947 ;
  assign n2681 = ~x960 & ~x963 ;
  assign n2682 = n2680 & n2681 ;
  assign n2683 = n2679 & n2682 ;
  assign n2663 = ~x614 & ~x616 ;
  assign n2664 = ~x642 & n2663 ;
  assign n2665 = x603 & n2664 ;
  assign n2666 = ~x661 & ~x662 ;
  assign n2667 = ~x681 & n2666 ;
  assign n2668 = x680 & n2667 ;
  assign n2669 = ~n2665 & ~n2668 ;
  assign n2684 = n2683 ^ n2669 ;
  assign n2685 = ~n2655 & n2684 ;
  assign n2686 = n2685 ^ n2683 ;
  assign n2687 = n2676 & ~n2686 ;
  assign n2656 = ~x969 & ~x971 ;
  assign n2657 = ~x974 & ~x977 ;
  assign n2658 = n2656 & n2657 ;
  assign n2659 = ~x587 & ~x602 ;
  assign n2660 = ~x961 & ~x967 ;
  assign n2661 = n2659 & n2660 ;
  assign n2662 = n2658 & n2661 ;
  assign n2670 = n2669 ^ n2662 ;
  assign n2671 = n2655 & n2670 ;
  assign n2672 = n2671 ^ n2669 ;
  assign n2673 = n1935 & ~n2672 ;
  assign n2688 = n2687 ^ n2673 ;
  assign n2689 = n2654 & n2688 ;
  assign n2693 = x829 & x1092 ;
  assign n2694 = ~n1847 & n2693 ;
  assign n2695 = ~n1849 & n2606 ;
  assign n2696 = n2695 ^ n2607 ;
  assign n2697 = ~n2694 & n2696 ;
  assign n2692 = n2608 ^ n1864 ;
  assign n2698 = n2697 ^ n2692 ;
  assign n2699 = ~x299 & n2655 ;
  assign n2700 = n2699 ^ n2655 ;
  assign n2701 = n2672 & ~n2700 ;
  assign n2702 = ~n2698 & n2701 ;
  assign n2703 = n2702 ^ n2698 ;
  assign n2704 = n2653 & ~n2703 ;
  assign n2705 = n1508 ^ n1419 ;
  assign n2706 = n2704 & ~n2705 ;
  assign n2707 = n2683 & n2700 ;
  assign n2708 = n2706 & ~n2707 ;
  assign n2711 = ~n2689 & ~n2708 ;
  assign n2712 = n2646 & n2711 ;
  assign n2713 = n2712 ^ n2646 ;
  assign n2714 = n2713 ^ n2645 ;
  assign n2715 = ~n1341 & ~n2714 ;
  assign n2716 = ~n2604 & ~n2715 ;
  assign n2732 = n2730 ^ n2716 ;
  assign n2742 = n2741 ^ n2732 ;
  assign n2769 = ~x58 & n1605 ;
  assign n2770 = ~x85 & n1716 ;
  assign n2771 = n1215 & n1680 ;
  assign n2772 = n1712 ^ n1210 ;
  assign n2775 = ~x67 & n2772 ;
  assign n2776 = n2775 ^ n1210 ;
  assign n2777 = n2771 & n2776 ;
  assign n2778 = ~n1678 & ~n2777 ;
  assign n2779 = n2770 & n2778 ;
  assign n2780 = ~x82 & ~n2721 ;
  assign n2781 = n2779 & n2780 ;
  assign n2782 = n2769 & ~n2781 ;
  assign n2762 = x103 & ~x109 ;
  assign n2763 = ~x314 & n2762 ;
  assign n2764 = n2763 ^ x109 ;
  assign n4884 = n1919 & n2764 ;
  assign n2759 = n1556 & n1746 ;
  assign n2760 = n1825 & n2759 ;
  assign n2761 = ~n1919 & ~n2760 ;
  assign n2786 = ~n4884 ^ n2761 ;
  assign n2787 = n2782 & n2786 ;
  assign n2788 = n2720 & n2787 ;
  assign n2789 = n2788 ^ n2720 ;
  assign n2767 = ~n4884 ^ n2720 ;
  assign n2790 = n2789 ^ n2767 ;
  assign n2791 = ~x72 & n2790 ;
  assign n2793 = n1265 & n1556 ;
  assign n2794 = n1611 & ~n1762 ;
  assign n2795 = n2793 & n2794 ;
  assign n2808 = n1265 & n1271 ;
  assign n2809 = x90 & n1561 ;
  assign n2810 = x841 & n2809 ;
  assign n2811 = n2810 ^ n1561 ;
  assign n2812 = n2808 & n2811 ;
  assign n2807 = ~n1786 & n2737 ;
  assign n2813 = n2812 ^ n2807 ;
  assign n2800 = ~x73 & n1269 ;
  assign n2801 = n1235 & n1238 ;
  assign n2802 = n1261 & n1639 ;
  assign n2803 = n2801 & n2802 ;
  assign n2804 = n2800 & n2803 ;
  assign n2805 = ~x32 & n1404 ;
  assign n2806 = n2804 & n2805 ;
  assign n2814 = n2813 ^ n2806 ;
  assign n2817 = ~n1272 & ~n2814 ;
  assign n2818 = n2795 & n2817 ;
  assign n2819 = n2818 ^ n2795 ;
  assign n2792 = n1556 & n1762 ;
  assign n2820 = n2819 ^ n2792 ;
  assign n2821 = ~n2791 & n2820 ;
  assign n2858 = ~x228 & n2821 ;
  assign n2859 = ~x228 & ~n1290 ;
  assign n2860 = n1340 & n2859 ;
  assign n2849 = ~x30 & x228 ;
  assign n2850 = ~n1290 & ~n2849 ;
  assign n2861 = n2860 ^ n2850 ;
  assign n2824 = n2653 & n2697 ;
  assign n2825 = n2674 ^ n1420 ;
  assign n2826 = n1281 & n2825 ;
  assign n2827 = n2824 & n2826 ;
  assign n2828 = n2827 ^ n1281 ;
  assign n2832 = n2676 ^ n1935 ;
  assign n2837 = n2828 & n2832 ;
  assign n2838 = n2654 & n2837 ;
  assign n2839 = n2838 ^ n2654 ;
  assign n2830 = n2827 ^ n2654 ;
  assign n2840 = n2839 ^ n2830 ;
  assign n2841 = n1273 & n2840 ;
  assign n2842 = ~x228 & ~n2841 ;
  assign n2843 = n1274 & n2635 ;
  assign n2844 = n1306 & n1328 ;
  assign n2845 = n1340 & n2844 ;
  assign n2846 = n2843 & n2845 ;
  assign n2847 = n2846 ^ n1340 ;
  assign n2848 = n2842 & n2847 ;
  assign n2851 = n2850 ^ n2849 ;
  assign n2852 = ~n2848 & ~n2851 ;
  assign n2862 = n2861 ^ n2852 ;
  assign n2863 = ~n2858 & ~n2862 ;
  assign n2872 = ~n2655 & n2668 ;
  assign n2864 = ~x299 & ~n2850 ;
  assign n2865 = x109 & ~x228 ;
  assign n2743 = x158 & x159 ;
  assign n2744 = x197 & n2743 ;
  assign n2745 = x160 & x232 ;
  assign n2746 = n2744 & n2745 ;
  assign n2866 = n2655 & n2746 ;
  assign n2867 = n2865 & n2866 ;
  assign n2868 = n2867 ^ n2655 ;
  assign n2869 = n2864 & n2868 ;
  assign n2870 = n2869 ^ n2868 ;
  assign n2871 = x907 & n2870 ;
  assign n2873 = n2872 ^ n2871 ;
  assign n2874 = ~n2863 & n2873 ;
  assign n2747 = x109 & x145 ;
  assign n2748 = x180 & x181 ;
  assign n2749 = n2747 & n2748 ;
  assign n2750 = x182 & x232 ;
  assign n2751 = n2749 & n2750 ;
  assign n2752 = n2751 ^ n2746 ;
  assign n2753 = x299 & n2752 ;
  assign n2754 = n2753 ^ n2751 ;
  assign n2755 = n2655 & n2754 ;
  assign n2756 = ~x109 & n2753 ;
  assign n2757 = n2755 & n2756 ;
  assign n2758 = n2757 ^ n2755 ;
  assign n2822 = ~n2758 & n2821 ;
  assign n2823 = ~x228 & n2822 ;
  assign n2854 = n2852 ^ n2823 ;
  assign n2855 = ~n2699 & n2854 ;
  assign n2856 = n2855 ^ n2854 ;
  assign n2857 = x602 & n2856 ;
  assign n2876 = n2874 ^ n2857 ;
  assign n2877 = n2665 ^ x947 ;
  assign n2878 = ~n2655 & n2877 ;
  assign n2879 = n2878 ^ x947 ;
  assign n2887 = ~n2855 & ~n2861 ;
  assign n2880 = n2879 ^ x587 ;
  assign n2881 = n2880 ^ n2855 ;
  assign n2882 = n2881 ^ n2854 ;
  assign n2888 = n2887 ^ n2882 ;
  assign n2889 = n2879 & n2888 ;
  assign n2890 = n2889 ^ n2882 ;
  assign n2891 = n2890 ^ x587 ;
  assign n2892 = n2890 ^ n2879 ;
  assign n2893 = ~n2889 & ~n2892 ;
  assign n2894 = ~n2891 & n2893 ;
  assign n2895 = n2894 ^ n2890 ;
  assign n2898 = x967 & n2856 ;
  assign n2896 = ~n2863 & n2870 ;
  assign n2897 = x970 & n2896 ;
  assign n2900 = n2898 ^ n2897 ;
  assign n2902 = x299 & x972 ;
  assign n2901 = ~x299 & x961 ;
  assign n2903 = n2902 ^ n2901 ;
  assign n2904 = n2902 ^ n2746 ;
  assign n2905 = n2904 ^ n2901 ;
  assign n2906 = n2905 ^ x109 ;
  assign n2916 = n2904 ^ n2752 ;
  assign n2917 = ~n2906 & n2916 ;
  assign n2918 = n2917 ^ n2902 ;
  assign n2920 = n2901 & n2916 ;
  assign n2921 = n2920 ^ n2905 ;
  assign n2922 = n2902 & ~n2921 ;
  assign n2923 = n2918 & n2922 ;
  assign n2924 = n2923 ^ n2920 ;
  assign n2925 = n2924 ^ n2746 ;
  assign n2926 = n2925 ^ n2905 ;
  assign n2927 = n2858 & n2926 ;
  assign n2928 = n2655 & ~n2927 ;
  assign n2929 = n2852 & n2928 ;
  assign n2930 = n2903 & n2929 ;
  assign n2931 = n2930 ^ n2928 ;
  assign n2933 = x972 & n2861 ;
  assign n2934 = n2931 & n2933 ;
  assign n2932 = n2931 ^ n2655 ;
  assign n2935 = n2934 ^ n2932 ;
  assign n2937 = x960 & n2896 ;
  assign n2936 = x977 & n2856 ;
  assign n2939 = n2937 ^ n2936 ;
  assign n2941 = x963 & n2896 ;
  assign n2940 = x969 & n2856 ;
  assign n2943 = n2941 ^ n2940 ;
  assign n2945 = x971 & n2856 ;
  assign n2944 = x975 & n2896 ;
  assign n2947 = n2945 ^ n2944 ;
  assign n2949 = x974 & n2856 ;
  assign n2948 = x978 & n2896 ;
  assign n2951 = n2949 ^ n2948 ;
  assign n2952 = ~x70 & n1261 ;
  assign n2953 = ~x96 & n1272 ;
  assign n2954 = n1268 & n2953 ;
  assign n2955 = n2952 & n2954 ;
  assign n2956 = n1244 & n2955 ;
  assign n2957 = ~x92 & n1450 ;
  assign n2958 = n1290 & n2957 ;
  assign n2959 = n2956 & n2958 ;
  assign n2960 = ~x39 & ~x72 ;
  assign n2961 = n2960 ^ x72 ;
  assign n2962 = n2959 & ~n2961 ;
  assign n2963 = x51 & ~x87 ;
  assign n2964 = n2963 ^ x87 ;
  assign n2965 = n1209 & ~n2964 ;
  assign n2966 = n2962 & n2965 ;
  assign n2973 = n1290 & n1420 ;
  assign n2974 = ~n2672 & n2973 ;
  assign n2971 = n1347 & ~n1537 ;
  assign n2972 = ~n2686 & n2971 ;
  assign n2975 = n2974 ^ n2972 ;
  assign n2976 = n2824 & n2975 ;
  assign n2981 = n2966 & ~n2976 ;
  assign n2982 = ~n2689 & n2981 ;
  assign n2983 = n2982 ^ n2689 ;
  assign n2968 = n2966 ^ n2847 ;
  assign n2969 = n2968 ^ n2689 ;
  assign n2984 = n2983 ^ n2969 ;
  assign n2985 = ~n2822 & n2984 ;
  assign n2986 = n2985 ^ x24 ;
  assign n2987 = ~x954 & n2986 ;
  assign n2988 = n2987 ^ x24 ;
  assign n2990 = n1303 & ~n1797 ;
  assign n2991 = n1499 & n2990 ;
  assign n2992 = n2991 ^ n1303 ;
  assign n2993 = n2992 ^ n1920 ;
  assign n2994 = n2993 ^ x105 ;
  assign n2995 = ~x228 & ~n2994 ;
  assign n2996 = n2995 ^ x105 ;
  assign n3000 = x119 & ~x468 ;
  assign n3001 = ~x1056 & n3000 ;
  assign n2997 = ~x119 & ~x228 ;
  assign n2998 = x252 & ~x468 ;
  assign n2999 = n2997 & n2998 ;
  assign n3002 = n3001 ^ n2999 ;
  assign n3003 = ~x1077 & n3000 ;
  assign n3004 = n3003 ^ n2999 ;
  assign n3005 = ~x1073 & n3000 ;
  assign n3006 = n3005 ^ n2999 ;
  assign n3007 = ~x1041 & n3000 ;
  assign n3008 = n3007 ^ n2999 ;
  assign n3013 = x1162 ^ x1161 ;
  assign n3010 = x1161 & x1162 ;
  assign n3014 = n3013 ^ n3010 ;
  assign n3015 = ~x590 & ~x592 ;
  assign n3021 = x390 ^ x324 ;
  assign n3022 = n3021 ^ x319 ;
  assign n3019 = x456 ^ x412 ;
  assign n3017 = x404 ^ x397 ;
  assign n3016 = x411 ^ x410 ;
  assign n3018 = n3017 ^ n3016 ;
  assign n3020 = n3019 ^ n3018 ;
  assign n3023 = n3022 ^ n3020 ;
  assign n3024 = x1196 & n3023 ;
  assign n3030 = x326 ^ x325 ;
  assign n3031 = n3030 ^ x318 ;
  assign n3028 = x405 ^ x403 ;
  assign n3026 = x409 ^ x406 ;
  assign n3025 = x402 ^ x401 ;
  assign n3027 = n3026 ^ n3025 ;
  assign n3029 = n3028 ^ n3027 ;
  assign n3032 = n3031 ^ n3029 ;
  assign n3033 = x1199 & n3032 ;
  assign n3034 = ~n3024 & ~n3033 ;
  assign n3035 = n3015 & ~n3034 ;
  assign n3041 = x421 ^ x420 ;
  assign n3042 = n3041 ^ x419 ;
  assign n3039 = x459 ^ x454 ;
  assign n3037 = x432 ^ x425 ;
  assign n3036 = x424 ^ x423 ;
  assign n3038 = n3037 ^ n3036 ;
  assign n3040 = n3039 ^ n3038 ;
  assign n3043 = n3042 ^ n3040 ;
  assign n3044 = x1198 & n3043 ;
  assign n3050 = x417 ^ x416 ;
  assign n3051 = n3050 ^ x415 ;
  assign n3048 = x464 ^ x453 ;
  assign n3046 = x431 ^ x418 ;
  assign n3045 = x438 ^ x437 ;
  assign n3047 = n3046 ^ n3045 ;
  assign n3049 = n3048 ^ n3047 ;
  assign n3052 = n3051 ^ n3049 ;
  assign n3053 = x1197 & n3052 ;
  assign n3054 = ~n3044 & ~n3053 ;
  assign n3060 = x428 ^ x427 ;
  assign n3061 = n3060 ^ x426 ;
  assign n3058 = x451 ^ x449 ;
  assign n3056 = x433 ^ x430 ;
  assign n3055 = x448 ^ x445 ;
  assign n3057 = n3056 ^ n3055 ;
  assign n3059 = n3058 ^ n3057 ;
  assign n3062 = n3061 ^ n3059 ;
  assign n3063 = x1199 & n3062 ;
  assign n3069 = x429 ^ x422 ;
  assign n3070 = n3069 ^ x414 ;
  assign n3067 = x443 ^ x436 ;
  assign n3065 = x446 ^ x444 ;
  assign n3064 = x435 ^ x434 ;
  assign n3066 = n3065 ^ n3064 ;
  assign n3068 = n3067 ^ n3066 ;
  assign n3071 = n3070 ^ n3068 ;
  assign n3072 = x1196 & n3071 ;
  assign n3073 = ~n3063 & ~n3072 ;
  assign n3074 = n3054 & n3073 ;
  assign n3075 = x588 & n3015 ;
  assign n3076 = ~n3074 & n3075 ;
  assign n3077 = n3076 ^ x588 ;
  assign n3079 = x591 & ~x592 ;
  assign n3078 = x592 ^ x590 ;
  assign n3080 = n3079 ^ n3078 ;
  assign n3126 = x353 ^ x352 ;
  assign n3127 = n3126 ^ x351 ;
  assign n3124 = x462 ^ x461 ;
  assign n3122 = x360 ^ x357 ;
  assign n3121 = x356 ^ x354 ;
  assign n3123 = n3122 ^ n3121 ;
  assign n3125 = n3124 ^ n3123 ;
  assign n3128 = n3127 ^ n3125 ;
  assign n3129 = x1199 & n3128 ;
  assign n3135 = x355 ^ x342 ;
  assign n3136 = n3135 ^ x320 ;
  assign n3133 = x455 ^ x452 ;
  assign n3131 = x460 ^ x458 ;
  assign n3130 = x441 ^ x361 ;
  assign n3132 = n3131 ^ n3130 ;
  assign n3134 = n3133 ^ n3132 ;
  assign n3137 = n3136 ^ n3134 ;
  assign n3138 = x1196 & n3137 ;
  assign n3139 = ~n3129 & ~n3138 ;
  assign n3145 = x321 ^ x316 ;
  assign n3146 = n3145 ^ x315 ;
  assign n3143 = x349 ^ x348 ;
  assign n3141 = x359 ^ x350 ;
  assign n3140 = x347 ^ x322 ;
  assign n3142 = n3141 ^ n3140 ;
  assign n3144 = n3143 ^ n3142 ;
  assign n3147 = n3146 ^ n3144 ;
  assign n3148 = x1198 & n3147 ;
  assign n3154 = x343 ^ x327 ;
  assign n3155 = n3154 ^ x323 ;
  assign n3152 = x450 ^ x362 ;
  assign n3150 = x358 ^ x346 ;
  assign n3149 = x345 ^ x344 ;
  assign n3151 = n3150 ^ n3149 ;
  assign n3153 = n3152 ^ n3151 ;
  assign n3156 = n3155 ^ n3153 ;
  assign n3157 = x1197 & n3156 ;
  assign n3158 = ~n3148 & ~n3157 ;
  assign n3159 = n3139 & n3158 ;
  assign n3086 = x371 ^ x370 ;
  assign n3087 = n3086 ^ x369 ;
  assign n3084 = x442 ^ x440 ;
  assign n3082 = x384 ^ x375 ;
  assign n3081 = x374 ^ x373 ;
  assign n3083 = n3082 ^ n3081 ;
  assign n3085 = n3084 ^ n3083 ;
  assign n3088 = n3087 ^ n3085 ;
  assign n3089 = x1198 & n3088 ;
  assign n3095 = x339 ^ x338 ;
  assign n3096 = n3095 ^ x337 ;
  assign n3093 = x388 ^ x387 ;
  assign n3091 = x372 ^ x363 ;
  assign n3090 = x386 ^ x380 ;
  assign n3092 = n3091 ^ n3090 ;
  assign n3094 = n3093 ^ n3092 ;
  assign n3097 = n3096 ^ n3094 ;
  assign n3098 = x1196 & n3097 ;
  assign n3099 = ~n3089 & ~n3098 ;
  assign n3105 = x365 ^ x364 ;
  assign n3106 = n3105 ^ x336 ;
  assign n3103 = x447 ^ x389 ;
  assign n3101 = x383 ^ x368 ;
  assign n3100 = x367 ^ x366 ;
  assign n3102 = n3101 ^ n3100 ;
  assign n3104 = n3103 ^ n3102 ;
  assign n3107 = n3106 ^ n3104 ;
  assign n3108 = x1197 & n3107 ;
  assign n3109 = n3099 & ~n3108 ;
  assign n3115 = x377 ^ x376 ;
  assign n3116 = n3115 ^ x317 ;
  assign n3113 = x382 ^ x381 ;
  assign n3111 = x439 ^ x385 ;
  assign n3110 = x379 ^ x378 ;
  assign n3112 = n3111 ^ n3110 ;
  assign n3114 = n3113 ^ n3112 ;
  assign n3117 = n3116 ^ n3114 ;
  assign n3118 = x1199 & n3117 ;
  assign n3119 = ~x591 & ~n3118 ;
  assign n3120 = n3109 & n3119 ;
  assign n3160 = n3159 ^ n3120 ;
  assign n9440 = ~x591 & ~x592 ;
  assign n3162 = n3160 & ~n9440 ;
  assign n3163 = n3162 ^ n3159 ;
  assign n3164 = n3080 & ~n3163 ;
  assign n3165 = ~n3077 & ~n3164 ;
  assign n3166 = n3165 ^ x588 ;
  assign n3167 = ~x217 & ~n3166 ;
  assign n3173 = x335 ^ x334 ;
  assign n3174 = n3173 ^ x333 ;
  assign n3171 = x463 ^ x413 ;
  assign n3169 = x407 ^ x393 ;
  assign n3168 = x392 ^ x391 ;
  assign n3170 = n3169 ^ n3168 ;
  assign n3172 = n3171 ^ n3170 ;
  assign n3175 = n3174 ^ n3172 ;
  assign n3176 = x1197 & n3175 ;
  assign n3182 = x394 ^ x329 ;
  assign n3183 = n3182 ^ x328 ;
  assign n3180 = x399 ^ x398 ;
  assign n3178 = x408 ^ x400 ;
  assign n3177 = x396 ^ x395 ;
  assign n3179 = n3178 ^ n3177 ;
  assign n3181 = n3180 ^ n3179 ;
  assign n3184 = n3183 ^ n3181 ;
  assign n3185 = x1198 & n3184 ;
  assign n3186 = ~n3176 & ~n3185 ;
  assign n3187 = n3079 & ~n3186 ;
  assign n3188 = n3187 ^ x591 ;
  assign n3189 = n3167 & n3188 ;
  assign n3190 = x567 & n3189 ;
  assign n3191 = n3035 & n3190 ;
  assign n3192 = n3191 ^ n3189 ;
  assign n3193 = n3192 ^ n3167 ;
  assign n3194 = ~n3014 & ~n3193 ;
  assign n3195 = ~x98 & x567 ;
  assign n3196 = ~x285 & ~x288 ;
  assign n3197 = ~x286 & ~x289 ;
  assign n3198 = n3196 & n3197 ;
  assign n3199 = n1847 & n2606 ;
  assign n3200 = ~x122 & n3199 ;
  assign n3201 = ~n3198 & n3200 ;
  assign n3202 = ~n1290 & n3201 ;
  assign n3203 = n3195 & n3202 ;
  assign n3204 = n3194 & n3203 ;
  assign n3009 = x1092 & x1093 ;
  assign n3011 = ~x31 & n3010 ;
  assign n3012 = n3009 & n3011 ;
  assign n3205 = n3204 ^ n3012 ;
  assign n3206 = ~x1163 & n3205 ;
  assign n3207 = n3009 & ~n3195 ;
  assign n3208 = n1290 & ~n3207 ;
  assign n3209 = ~x1163 & ~n3014 ;
  assign n3260 = x100 ^ x39 ;
  assign n3263 = ~x35 & ~x70 ;
  assign n3264 = x90 ^ x51 ;
  assign n3265 = n3264 ^ x93 ;
  assign n3266 = x93 ^ x90 ;
  assign n3267 = x841 ^ x93 ;
  assign n3270 = n3266 & ~n3267 ;
  assign n3271 = n3270 ^ x90 ;
  assign n3272 = n3265 & ~n3271 ;
  assign n3273 = n3263 & n3272 ;
  assign n3274 = n1262 & n3273 ;
  assign n3261 = n1264 & n1745 ;
  assign n3262 = x98 & n3261 ;
  assign n3276 = n3274 ^ n3262 ;
  assign n3277 = ~x96 & ~n3276 ;
  assign n3278 = ~x72 & n2608 ;
  assign n3286 = ~x98 & n3278 ;
  assign n3287 = x1091 & n3286 ;
  assign n3288 = n3287 ^ x1091 ;
  assign n3279 = n3278 ^ x72 ;
  assign n3280 = n3279 ^ x1091 ;
  assign n3289 = n3288 ^ n3280 ;
  assign n3290 = ~n2698 & ~n3289 ;
  assign n3291 = ~n3277 & n3290 ;
  assign n3292 = x91 & n1810 ;
  assign n3293 = ~x24 & ~x58 ;
  assign n3294 = n3292 & n3293 ;
  assign n3295 = n3294 ^ n1857 ;
  assign n3296 = ~x72 & n1264 ;
  assign n3218 = ~x122 & n1864 ;
  assign n3297 = n1268 & n3218 ;
  assign n3298 = n3296 & n3297 ;
  assign n3299 = n3295 & n3298 ;
  assign n3300 = ~n3291 & ~n3299 ;
  assign n3301 = n1264 & n1752 ;
  assign n3302 = ~x122 & x829 ;
  assign n3303 = ~x841 & n1272 ;
  assign n3304 = n3302 & n3303 ;
  assign n3305 = n3301 & n3304 ;
  assign n3306 = ~n2953 & ~n3305 ;
  assign n3307 = ~n3300 & ~n3306 ;
  assign n3308 = ~x75 & ~n3307 ;
  assign n3309 = ~n3260 & n3308 ;
  assign n3317 = n2953 & n2960 ;
  assign n3318 = ~x87 & n3276 ;
  assign n3319 = n3317 & n3318 ;
  assign n3320 = n3319 ^ x87 ;
  assign n3325 = ~n2698 & n3320 ;
  assign n3247 = ~x87 & n3218 ;
  assign n3248 = ~x24 & ~x100 ;
  assign n3219 = x232 & n2655 ;
  assign n3220 = n1793 & ~n2619 ;
  assign n3221 = n3219 & n3220 ;
  assign n3222 = n3221 ^ n2619 ;
  assign n3249 = x252 & n3222 ;
  assign n3250 = n3249 ^ x252 ;
  assign n3251 = n3248 & n3250 ;
  assign n3252 = n3247 & n3251 ;
  assign n3253 = n1273 & n3252 ;
  assign n3254 = x75 & ~n3253 ;
  assign n3255 = ~x39 & ~x100 ;
  assign n3256 = n1273 & n1279 ;
  assign n3257 = n3255 & n3256 ;
  assign n3258 = ~n3254 & n3257 ;
  assign n3311 = n3309 ^ n3258 ;
  assign n3210 = ~x87 & ~x92 ;
  assign n3211 = n3210 ^ x100 ;
  assign n3212 = n1293 & ~n3211 ;
  assign n3223 = n3218 & ~n3222 ;
  assign n3226 = n3212 & n3223 ;
  assign n3227 = x228 & n3226 ;
  assign n3228 = n3227 ^ x228 ;
  assign n3213 = n3212 ^ n1293 ;
  assign n3214 = n3213 ^ x228 ;
  assign n3229 = n3228 ^ n3214 ;
  assign n3230 = n3210 & n3229 ;
  assign n3231 = n1273 & n3230 ;
  assign n3232 = n3231 ^ x39 ;
  assign n3233 = n2675 ^ n1421 ;
  assign n3236 = n1510 & ~n2686 ;
  assign n3234 = n1423 & ~n2672 ;
  assign n3237 = n3236 ^ n3234 ;
  assign n3238 = n3233 & n3237 ;
  assign n3239 = n2654 & n3238 ;
  assign n3240 = n3239 ^ n1280 ;
  assign n3243 = n3231 & ~n3240 ;
  assign n3244 = n3243 ^ n1280 ;
  assign n3245 = ~n3232 & ~n3244 ;
  assign n3246 = n3245 ^ x39 ;
  assign n3312 = n3311 ^ n3246 ;
  assign n3326 = n3325 ^ n3312 ;
  assign n3327 = n3309 & ~n3326 ;
  assign n3328 = n3327 ^ n3312 ;
  assign n3329 = n3328 ^ n3309 ;
  assign n3330 = n3309 ^ n3246 ;
  assign n3331 = ~n3327 & ~n3330 ;
  assign n3332 = n3329 & n3331 ;
  assign n3333 = n3332 ^ n3328 ;
  assign n3334 = n1847 & n3193 ;
  assign n3335 = ~n3333 & n3334 ;
  assign n3336 = n3335 ^ n3333 ;
  assign n3337 = ~n3198 & n3336 ;
  assign n3345 = ~n3188 & n3337 ;
  assign n3346 = n3167 & n3345 ;
  assign n3347 = n3346 ^ n3167 ;
  assign n3338 = n3337 ^ n3336 ;
  assign n3339 = n3338 ^ n3167 ;
  assign n3348 = n3347 ^ n3339 ;
  assign n3349 = n3209 & ~n3348 ;
  assign n3350 = n3208 & n3349 ;
  assign n3358 = ~x217 & ~x588 ;
  assign n3359 = x591 & ~x1091 ;
  assign n3360 = n3358 & n3359 ;
  assign n3361 = n3186 & n3360 ;
  assign n3362 = n3035 & n3361 ;
  assign n3355 = x567 & n2608 ;
  assign n3351 = n3199 & n3317 ;
  assign n3352 = n3351 ^ n3260 ;
  assign n3353 = n3274 & n3352 ;
  assign n3354 = n3353 ^ n3260 ;
  assign n3356 = n3355 ^ n3354 ;
  assign n3357 = n3356 ^ n3307 ;
  assign n3363 = n3362 ^ n3355 ;
  assign n3364 = n3363 ^ n3307 ;
  assign n3365 = n3362 ^ x1199 ;
  assign n3366 = n3365 ^ n3354 ;
  assign n3367 = n3364 & ~n3366 ;
  assign n3368 = n3357 & n3367 ;
  assign n3369 = n3368 ^ n3362 ;
  assign n3370 = n3369 ^ n3354 ;
  assign n3371 = ~n3307 & n3370 ;
  assign n3372 = n3354 & n3371 ;
  assign n3373 = n3372 ^ n3307 ;
  assign n3374 = ~n3246 & n3373 ;
  assign n3411 = n3200 ^ n2698 ;
  assign n3376 = n3200 ^ x98 ;
  assign n3412 = n3411 ^ n3376 ;
  assign n3415 = n3412 ^ n1276 ;
  assign n3413 = n3412 ^ n3258 ;
  assign n3414 = n3413 ^ n3376 ;
  assign n3433 = n3415 ^ n3414 ;
  assign n3434 = n3433 ^ n3411 ;
  assign n3435 = n3434 ^ n3200 ;
  assign n3416 = n3415 ^ n3376 ;
  assign n3417 = n3416 ^ n3414 ;
  assign n3394 = ~n3200 & ~n3376 ;
  assign n3395 = n3413 ^ n3394 ;
  assign n3396 = n3412 ^ n3395 ;
  assign n3397 = n3396 ^ x98 ;
  assign n3399 = n3434 ^ x98 ;
  assign n3400 = ~n3397 & n3399 ;
  assign n3385 = n3433 ^ n3412 ;
  assign n3401 = n3415 ^ n3385 ;
  assign n3402 = n3435 ^ n3401 ;
  assign n3403 = n3413 ^ n3385 ;
  assign n3404 = n3435 ^ n3403 ;
  assign n3405 = ~n3402 & n3404 ;
  assign n3406 = n3400 & n3405 ;
  assign n3407 = n3406 ^ n3394 ;
  assign n3408 = n3417 ^ n3407 ;
  assign n3429 = n3408 ^ n2698 ;
  assign n3430 = n3435 ^ n3429 ;
  assign n3431 = n3430 ^ n3417 ;
  assign n3438 = n3431 ^ n2698 ;
  assign n3439 = n3438 ^ x98 ;
  assign n3440 = n3439 ^ n3435 ;
  assign n3441 = ~n3374 & ~n3440 ;
  assign n3449 = n3355 & n3441 ;
  assign n3450 = n3362 & n3449 ;
  assign n3451 = n3450 ^ n3362 ;
  assign n3442 = n3441 ^ n3374 ;
  assign n3443 = n3442 ^ n3362 ;
  assign n3452 = n3451 ^ n3443 ;
  assign n3453 = n3350 & n3452 ;
  assign n3454 = ~n3206 & ~n3453 ;
  assign n3455 = x76 & ~n1728 ;
  assign n3459 = ~x137 & ~n1784 ;
  assign n3462 = ~n1851 & ~n3198 ;
  assign n3465 = n3459 & ~n3462 ;
  assign n3466 = n3455 & n3465 ;
  assign n3467 = n3466 ^ n3455 ;
  assign n3456 = ~x24 & n1245 ;
  assign n3457 = n3456 ^ n3455 ;
  assign n3468 = n3467 ^ n3457 ;
  assign n3469 = ~x50 & n3468 ;
  assign n3470 = n3469 ^ n3456 ;
  assign n3471 = ~n1785 & ~n3470 ;
  assign n3474 = x32 & ~x841 ;
  assign n3477 = ~x24 & n3474 ;
  assign n3478 = n3477 ^ x32 ;
  assign n3479 = n3471 & n3478 ;
  assign n3480 = n3479 ^ n3470 ;
  assign n3481 = n1919 & n3480 ;
  assign n3491 = x75 & n3248 ;
  assign n3492 = n1851 & n3491 ;
  assign n3493 = n3492 ^ n3491 ;
  assign n3496 = n3222 & n3493 ;
  assign n3483 = n2608 ^ x129 ;
  assign n3484 = n2605 & n3483 ;
  assign n3485 = n3484 ^ x129 ;
  assign n3486 = n1274 & n3485 ;
  assign n3490 = ~n1797 & n3486 ;
  assign n3497 = n3496 ^ n3490 ;
  assign n3498 = x252 & n3497 ;
  assign n3499 = n3498 ^ n3490 ;
  assign n3494 = n3493 ^ n3486 ;
  assign n3500 = n3499 ^ n3494 ;
  assign n3501 = ~x137 & ~n3222 ;
  assign n3509 = ~n1797 & n3501 ;
  assign n3510 = n3493 & n3509 ;
  assign n3511 = n3510 ^ n3493 ;
  assign n3502 = n3501 ^ x137 ;
  assign n3503 = n3502 ^ n3493 ;
  assign n3512 = n3511 ^ n3503 ;
  assign n3513 = n3500 & ~n3512 ;
  assign n3514 = n2844 & n3513 ;
  assign n3515 = ~n3481 & ~n3514 ;
  assign n3531 = x186 ^ x164 ;
  assign n3532 = ~x299 & n3531 ;
  assign n3533 = n3532 ^ x164 ;
  assign n3534 = ~n1277 & n3219 ;
  assign n3535 = n3533 & n3534 ;
  assign n3536 = n3535 ^ n1277 ;
  assign n3537 = n1271 & n2804 ;
  assign n3538 = n1310 & n3537 ;
  assign n3539 = ~x63 & ~x107 ;
  assign n3540 = ~x40 & n3539 ;
  assign n3557 = x176 ^ x154 ;
  assign n3560 = x299 & n3557 ;
  assign n3561 = n3560 ^ x176 ;
  assign n3562 = n3219 & n3561 ;
  assign n3567 = x92 & n3562 ;
  assign n3568 = n3540 & n3567 ;
  assign n3569 = n3568 ^ n3540 ;
  assign n3550 = x954 ^ x33 ;
  assign n3541 = ~x79 & ~x118 ;
  assign n3542 = ~x33 & ~x34 ;
  assign n3543 = n3541 & n3542 ;
  assign n3544 = ~x954 & n3543 ;
  assign n3545 = ~x138 & x139 ;
  assign n3546 = n3545 ^ x138 ;
  assign n3547 = n3544 & ~n3546 ;
  assign n3548 = ~x196 & n3547 ;
  assign n3549 = ~x195 & n3548 ;
  assign n3551 = n3550 ^ n3549 ;
  assign n3552 = n3540 & n3551 ;
  assign n3553 = ~x39 & n3210 ;
  assign n3554 = n3552 & ~n3553 ;
  assign n3555 = n3554 ^ n3540 ;
  assign n3570 = n3569 ^ n3555 ;
  assign n3571 = n3538 & n3570 ;
  assign n3572 = n3571 ^ n3554 ;
  assign n3573 = n3210 & n3301 ;
  assign n3574 = n3317 & n3573 ;
  assign n3575 = x38 & ~n3574 ;
  assign n3576 = ~x54 & ~n3575 ;
  assign n3577 = n3572 & n3576 ;
  assign n3581 = x39 & n3219 ;
  assign n3582 = n3219 ^ n1273 ;
  assign n3585 = n2676 & ~n2683 ;
  assign n3586 = ~x152 & n3585 ;
  assign n3583 = n1935 & ~n2662 ;
  assign n3584 = ~x174 & n3583 ;
  assign n3587 = n3586 ^ n3584 ;
  assign n3588 = n2824 & n3587 ;
  assign n3590 = x154 & n3585 ;
  assign n3589 = x176 & n3583 ;
  assign n3591 = n3590 ^ n3589 ;
  assign n3592 = n2654 & n3591 ;
  assign n3593 = ~n3588 & ~n3592 ;
  assign n3594 = n3593 ^ n3581 ;
  assign n3595 = ~n3582 & n3594 ;
  assign n3596 = n3581 & ~n3595 ;
  assign n3597 = n3596 ^ n3219 ;
  assign n3600 = n2824 ^ n2654 ;
  assign n3601 = n2688 & n3600 ;
  assign n3602 = n3537 & n3601 ;
  assign n3603 = n3210 & n3602 ;
  assign n3606 = ~n3597 & n3603 ;
  assign n3607 = n3577 & n3606 ;
  assign n3608 = n3607 ^ n3577 ;
  assign n3609 = n3608 ^ n3576 ;
  assign n3610 = n3536 & ~n3609 ;
  assign n3524 = x191 ^ x169 ;
  assign n3527 = x299 & n3524 ;
  assign n3528 = n3527 ^ x191 ;
  assign n3529 = n3219 & n3528 ;
  assign n3611 = n3610 ^ n3529 ;
  assign n3612 = ~x74 & n3611 ;
  assign n3517 = x183 ^ x178 ;
  assign n3516 = x157 ^ x149 ;
  assign n3518 = n3517 ^ n3516 ;
  assign n3521 = ~x299 & n3518 ;
  assign n3522 = n3521 ^ n3516 ;
  assign n3523 = n3219 & n3522 ;
  assign n3530 = n3529 ^ n3523 ;
  assign n3613 = n3612 ^ n3530 ;
  assign n3614 = ~n1275 & ~n3613 ;
  assign n3615 = n3614 ^ n3523 ;
  assign n3616 = n1290 & n3615 ;
  assign n3617 = n1314 & n3536 ;
  assign n3618 = x73 & n2803 ;
  assign n3619 = n1269 & n1271 ;
  assign n3620 = n3618 & n3619 ;
  assign n3623 = n1611 & n2814 ;
  assign n3621 = ~x70 & n1582 ;
  assign n3622 = n1762 & ~n3621 ;
  assign n3625 = n3623 ^ n3622 ;
  assign n3626 = ~n3620 & ~n3625 ;
  assign n3627 = n3552 & n3626 ;
  assign n3628 = n3617 & n3627 ;
  assign n3629 = n3616 & ~n3628 ;
  assign n3630 = n1280 & n3597 ;
  assign n3631 = n1611 & n2812 ;
  assign n3632 = x193 ^ x172 ;
  assign n3635 = x299 & n3632 ;
  assign n3636 = n3635 ^ x193 ;
  assign n3637 = n3631 & n3636 ;
  assign n3643 = ~x210 & n3474 ;
  assign n3644 = n3621 & n3643 ;
  assign n3645 = n3644 ^ n3621 ;
  assign n3650 = x149 & ~n3645 ;
  assign n3651 = x299 & n3650 ;
  assign n3652 = n3651 ^ x299 ;
  assign n3638 = x174 ^ x152 ;
  assign n3639 = ~x299 & n3638 ;
  assign n3640 = n3639 ^ x152 ;
  assign n3641 = n3640 ^ x299 ;
  assign n3653 = n3652 ^ n3641 ;
  assign n3654 = ~x73 & ~n3653 ;
  assign n3655 = n3654 ^ n3640 ;
  assign n3656 = x180 ^ x158 ;
  assign n3657 = ~x299 & n3656 ;
  assign n3658 = n3657 ^ x158 ;
  assign n3659 = n1270 & n3658 ;
  assign n3660 = n1404 & n3659 ;
  assign n3661 = n3660 ^ n3655 ;
  assign n3662 = n3655 & n3661 ;
  assign n3663 = ~n3637 & n3662 ;
  assign n3664 = n1774 & n3663 ;
  assign n3668 = ~x198 & ~x841 ;
  assign n1780 = n1271 ^ x95 ;
  assign n3669 = ~n1780 & n2804 ;
  assign n3670 = n3668 & n3669 ;
  assign n3671 = ~x299 & n3621 ;
  assign n3672 = ~n3670 & n3671 ;
  assign n3673 = n3672 ^ x299 ;
  assign n3678 = n3664 & ~n3673 ;
  assign n3679 = x183 & n3678 ;
  assign n3680 = n3679 ^ x183 ;
  assign n3665 = n3664 ^ n1774 ;
  assign n3666 = n3665 ^ x183 ;
  assign n3681 = n3680 ^ n3666 ;
  assign n3682 = ~x39 & ~n3681 ;
  assign n3683 = n3630 & ~n3682 ;
  assign n3684 = n3629 & ~n3683 ;
  assign n3687 = ~n1206 & n1277 ;
  assign n3692 = x164 & ~n3687 ;
  assign n3693 = n3692 ^ x169 ;
  assign n3694 = ~x74 & n3693 ;
  assign n3685 = n3516 ^ x169 ;
  assign n3695 = n3694 ^ n3685 ;
  assign n3696 = ~n1275 & n3695 ;
  assign n3697 = n3696 ^ n3516 ;
  assign n3698 = n3219 & n3697 ;
  assign n3699 = n3698 ^ n1275 ;
  assign n3700 = ~n1290 & ~n3699 ;
  assign n3701 = n1448 & ~n3687 ;
  assign n3702 = n3701 ^ n1448 ;
  assign n3703 = n3540 & n3702 ;
  assign n3706 = x149 & n3219 ;
  assign n3707 = n3706 ^ n3551 ;
  assign n3708 = n1325 & n3707 ;
  assign n3709 = n3708 ^ n3551 ;
  assign n3710 = n3703 & n3709 ;
  assign n3711 = n3700 & ~n3710 ;
  assign n3712 = ~n3684 & ~n3711 ;
  assign n3713 = ~x33 & ~x954 ;
  assign n3714 = n3713 ^ x34 ;
  assign n3715 = n3714 ^ n3549 ;
  assign n3717 = n1288 & n3537 ;
  assign n3718 = n3553 & n3717 ;
  assign n3719 = ~n1289 & ~n3718 ;
  assign n3716 = n1556 & n3626 ;
  assign n3720 = n3719 ^ n3716 ;
  assign n3721 = ~n3715 & n3720 ;
  assign n3723 = ~x161 & n3585 ;
  assign n3722 = ~x144 & n3583 ;
  assign n3724 = n3723 ^ n3722 ;
  assign n3725 = n2697 & n3724 ;
  assign n3727 = x155 & n3585 ;
  assign n3726 = x177 & n3583 ;
  assign n3728 = n3727 ^ n3726 ;
  assign n3729 = n1864 & n3728 ;
  assign n3730 = ~n3725 & ~n3729 ;
  assign n3731 = n3219 & ~n3730 ;
  assign n3732 = n3603 & ~n3731 ;
  assign n3733 = ~n1282 & n1289 ;
  assign n3734 = ~n3732 & n3733 ;
  assign n3735 = x92 & n3538 ;
  assign n3738 = x177 ^ x155 ;
  assign n3739 = ~x299 & n3738 ;
  assign n3740 = n3739 ^ x155 ;
  assign n3741 = n3219 & n3740 ;
  assign n3742 = n3741 ^ n3715 ;
  assign n3743 = n3735 & ~n3742 ;
  assign n3744 = n3743 ^ n3715 ;
  assign n3745 = n3734 & ~n3744 ;
  assign n3746 = n3745 ^ n3734 ;
  assign n3754 = n3603 & n3746 ;
  assign n3755 = x39 & n3754 ;
  assign n3756 = n3755 ^ x39 ;
  assign n3748 = n3745 ^ x39 ;
  assign n3757 = n3756 ^ n3748 ;
  assign n3758 = ~n3721 & ~n3757 ;
  assign n3759 = n3703 & ~n3758 ;
  assign n3788 = x145 ^ x140 ;
  assign n3786 = ~x178 & ~x183 ;
  assign n3784 = x197 ^ x162 ;
  assign n3783 = ~x149 & ~x157 ;
  assign n3785 = n3784 ^ n3783 ;
  assign n3787 = n3786 ^ n3785 ;
  assign n3789 = n3788 ^ n3787 ;
  assign n3790 = n1537 & n3789 ;
  assign n3791 = n3790 ^ n3785 ;
  assign n3766 = x148 ^ x141 ;
  assign n3767 = x299 & n3766 ;
  assign n3768 = n3767 ^ x141 ;
  assign n3760 = x188 ^ x167 ;
  assign n3763 = x299 & n3760 ;
  assign n3764 = n3763 ^ x188 ;
  assign n3765 = ~n3576 & n3764 ;
  assign n3769 = n3768 ^ n3765 ;
  assign n3770 = ~x74 & n3769 ;
  assign n3771 = n3770 ^ n3768 ;
  assign n3792 = n3791 ^ n3771 ;
  assign n3778 = x167 & ~n3687 ;
  assign n3779 = n3778 ^ x148 ;
  assign n3780 = ~x74 & n3779 ;
  assign n3772 = n3771 ^ x148 ;
  assign n3781 = n3780 ^ n3772 ;
  assign n3782 = ~n1290 & n3781 ;
  assign n3793 = n3792 ^ n3782 ;
  assign n3794 = ~n1275 & ~n3793 ;
  assign n3795 = n3794 ^ n3791 ;
  assign n3804 = x162 & x299 ;
  assign n3796 = x161 ^ x144 ;
  assign n3801 = x299 & n3796 ;
  assign n3802 = n3801 ^ x144 ;
  assign n3803 = x73 & ~n3802 ;
  assign n3805 = ~n3645 & ~n3803 ;
  assign n3806 = n3804 & n3805 ;
  assign n3807 = n3806 ^ n3803 ;
  assign n3808 = x181 ^ x159 ;
  assign n3809 = ~x299 & n3808 ;
  assign n3810 = n3809 ^ x159 ;
  assign n3811 = n2805 & n3810 ;
  assign n3812 = ~n3807 & n3811 ;
  assign n3813 = n3812 ^ x140 ;
  assign n3814 = n3812 ^ n3807 ;
  assign n3815 = n1919 & ~n3814 ;
  assign n3816 = ~n3673 & n3815 ;
  assign n3817 = n3813 & n3816 ;
  assign n3818 = n3817 ^ n3815 ;
  assign n3826 = ~n1796 & n3818 ;
  assign n3827 = n3631 & n3826 ;
  assign n3828 = n3827 ^ n3631 ;
  assign n3819 = n3818 ^ n1919 ;
  assign n3820 = n3819 ^ n3631 ;
  assign n3829 = n3828 ^ n3820 ;
  assign n3830 = n3795 & ~n3829 ;
  assign n3831 = n3219 & n3830 ;
  assign n3835 = n1342 & n3718 ;
  assign n3840 = n3831 & n3835 ;
  assign n3841 = x162 & n3840 ;
  assign n3842 = n3841 ^ x162 ;
  assign n3832 = n3831 ^ n3219 ;
  assign n3833 = n3832 ^ x162 ;
  assign n3843 = n3842 ^ n3833 ;
  assign n3844 = ~n3759 & ~n3843 ;
  assign n3881 = n1314 & ~n3574 ;
  assign n3882 = ~n3687 & n3881 ;
  assign n3883 = n3882 ^ n1313 ;
  assign n3857 = n1277 & n3486 ;
  assign n3845 = n1797 & ~n2619 ;
  assign n3860 = x683 & n2695 ;
  assign n3861 = n3860 ^ x137 ;
  assign n3862 = ~n3222 & n3861 ;
  assign n3863 = n3862 ^ x137 ;
  assign n3864 = x252 & n3863 ;
  assign n3865 = n3864 ^ x252 ;
  assign n3866 = ~n3845 & ~n3865 ;
  assign n3867 = n3857 & n3866 ;
  assign n3876 = n1797 & n3867 ;
  assign n3877 = ~x137 & n3876 ;
  assign n3878 = n3877 ^ x137 ;
  assign n3846 = x75 ^ x38 ;
  assign n3847 = n3846 ^ n3249 ;
  assign n3848 = ~n3845 & n3847 ;
  assign n3850 = x137 & ~n1851 ;
  assign n3851 = n3848 & n3850 ;
  assign n3849 = n3848 ^ n3845 ;
  assign n3852 = n3851 ^ n3849 ;
  assign n3853 = x75 & n3846 ;
  assign n3854 = n3852 & n3853 ;
  assign n3855 = n3854 ^ n3846 ;
  assign n3856 = n3248 & n3855 ;
  assign n3869 = n3867 ^ n3856 ;
  assign n3870 = n3869 ^ x137 ;
  assign n3879 = n3878 ^ n3870 ;
  assign n3880 = n3574 & n3879 ;
  assign n3884 = n3883 ^ n3880 ;
  assign n3885 = x24 & ~x59 ;
  assign n3886 = x40 & x1082 ;
  assign n3888 = ~x122 & n2608 ;
  assign n3889 = ~n3462 & n3888 ;
  assign n3890 = ~n3459 & n3889 ;
  assign n3891 = x76 & n3890 ;
  assign n3892 = n3891 ^ n1810 ;
  assign n3893 = n2782 & n3892 ;
  assign n3901 = n3267 & n3893 ;
  assign n3902 = n1558 & n3901 ;
  assign n3903 = n3902 ^ n1558 ;
  assign n3894 = n3893 ^ n3892 ;
  assign n3895 = n3894 ^ n1558 ;
  assign n3904 = n3903 ^ n3895 ;
  assign n3905 = ~n3886 & ~n3904 ;
  assign n3906 = n1774 & ~n3905 ;
  assign n3907 = ~n3885 & ~n3906 ;
  assign n3915 = ~n2807 & n3907 ;
  assign n3916 = n1318 & n3915 ;
  assign n3917 = n3916 ^ n1318 ;
  assign n3908 = n3907 ^ n3906 ;
  assign n3909 = n3908 ^ n1318 ;
  assign n3918 = n3917 ^ n3909 ;
  assign n3919 = n3884 & ~n3918 ;
  assign n3920 = n3919 ^ n3883 ;
  assign n3921 = ~x55 & ~x74 ;
  assign n3922 = n3885 ^ x24 ;
  assign n3923 = n1320 & ~n3922 ;
  assign n3924 = n3921 & n3923 ;
  assign n3925 = n3920 & n3924 ;
  assign n3926 = x36 & n1261 ;
  assign n3927 = ~n1728 & n3926 ;
  assign n3928 = ~n3294 & ~n3927 ;
  assign n3929 = n1268 & n2759 ;
  assign n3930 = ~n2608 & n3929 ;
  assign n3931 = ~n3928 & n3930 ;
  assign n3932 = ~x70 & ~x89 ;
  assign n3933 = x332 & n3932 ;
  assign n3934 = n3933 ^ x332 ;
  assign n3935 = n1261 & n3929 ;
  assign n3936 = ~n1728 & n3935 ;
  assign n3937 = x841 & n3936 ;
  assign n3938 = n3937 ^ n3936 ;
  assign n3947 = n3934 & n3938 ;
  assign n3939 = n1651 & n3935 ;
  assign n3940 = x64 & n3939 ;
  assign n3941 = x841 & n3940 ;
  assign n3942 = n3941 ^ n3940 ;
  assign n3943 = ~x24 & n1309 ;
  assign n3944 = n3943 ^ n1309 ;
  assign n3945 = ~n3942 & ~n3944 ;
  assign n3948 = n3947 ^ n3945 ;
  assign n3984 = n1785 & n2737 ;
  assign n3985 = n1556 & n3984 ;
  assign n3949 = ~x35 & ~x48 ;
  assign n3950 = ~x986 & n2608 ;
  assign n3951 = x252 & ~n3950 ;
  assign n3952 = x108 & x314 ;
  assign n3953 = ~n3951 & n3952 ;
  assign n3958 = ~x47 & ~n3953 ;
  assign n3959 = n3958 ^ x841 ;
  assign n3960 = n3949 & n3959 ;
  assign n3961 = n3960 ^ x841 ;
  assign n3962 = n2792 & ~n3961 ;
  assign n3963 = x287 & n2965 ;
  assign n3964 = n2962 & n3963 ;
  assign n3965 = n3964 ^ n2966 ;
  assign n3966 = x835 & ~x979 ;
  assign n3967 = x984 & n3966 ;
  assign n3968 = n3967 ^ x979 ;
  assign n3969 = n2651 & ~n3968 ;
  assign n3970 = n3969 ^ n3968 ;
  assign n3971 = x835 & ~n2703 ;
  assign n3972 = ~n2707 & n3971 ;
  assign n3977 = ~x1093 & ~n2706 ;
  assign n3973 = x786 & ~x1082 ;
  assign n3974 = ~n3970 & n3973 ;
  assign n3978 = n3977 ^ n3974 ;
  assign n3979 = n3972 & ~n3978 ;
  assign n3980 = n3979 ^ n3974 ;
  assign n3981 = ~n3970 & ~n3980 ;
  assign n3982 = n3965 & n3981 ;
  assign n3983 = ~n3962 & ~n3982 ;
  assign n3987 = n3985 ^ n3983 ;
  assign n3988 = x102 ^ x40 ;
  assign n3989 = n1919 & ~n3886 ;
  assign n3990 = n3988 & n3989 ;
  assign n4042 = n2959 & n3219 ;
  assign n4043 = n3963 & n4042 ;
  assign n4044 = n4043 ^ n3219 ;
  assign n4045 = ~n2961 & n4044 ;
  assign n4047 = ~x166 & ~n1537 ;
  assign n4049 = x152 & n4047 ;
  assign n4046 = n1483 & ~n1537 ;
  assign n4048 = n4047 ^ n4046 ;
  assign n4050 = n4049 ^ n4048 ;
  assign n4051 = n4050 ^ n4044 ;
  assign n4054 = ~x189 & n1537 ;
  assign n4056 = x174 & n4054 ;
  assign n4052 = n1468 & n1537 ;
  assign n4053 = n4052 ^ n4045 ;
  assign n4055 = n4054 ^ n4053 ;
  assign n4057 = n4056 ^ n4055 ;
  assign n4058 = n4051 & n4057 ;
  assign n4059 = n4045 & ~n4058 ;
  assign n4060 = n4059 ^ n2961 ;
  assign n3991 = n1279 & n1290 ;
  assign n3992 = x100 ^ x87 ;
  assign n3993 = n1273 ^ x87 ;
  assign n3994 = n3992 & ~n3993 ;
  assign n3995 = n3994 ^ x87 ;
  assign n3996 = n3991 & ~n3995 ;
  assign n3997 = ~n3254 & n3996 ;
  assign n3998 = ~n3306 & n3997 ;
  assign n3999 = n3261 ^ x228 ;
  assign n4000 = x110 ^ x94 ;
  assign n4002 = ~x250 & x252 ;
  assign n4003 = x901 & ~x959 ;
  assign n4004 = n4002 & n4003 ;
  assign n4001 = ~x480 & x949 ;
  assign n4005 = n4004 ^ n4001 ;
  assign n4006 = x110 & n4005 ;
  assign n4007 = n4006 ^ n4004 ;
  assign n4008 = n4000 & n4007 ;
  assign n4011 = n3999 & ~n4008 ;
  assign n4012 = n4011 ^ n3261 ;
  assign n4013 = n3998 & n4012 ;
  assign n4014 = x228 & ~n3299 ;
  assign n4019 = n1274 & ~n3223 ;
  assign n4020 = n4019 ^ n1276 ;
  assign n4021 = n4014 & n4020 ;
  assign n4022 = ~n3277 & n4021 ;
  assign n4029 = ~n1263 & ~n1851 ;
  assign n4030 = n4022 & n4029 ;
  assign n4031 = n4030 ^ n4022 ;
  assign n4032 = n4031 ^ n4021 ;
  assign n4033 = n4013 & ~n4032 ;
  assign n4034 = ~x44 & n4033 ;
  assign n4039 = ~x101 & n4034 ;
  assign n4040 = n4039 ^ x41 ;
  assign n4041 = n2960 & ~n4040 ;
  assign n4061 = n4060 ^ n4041 ;
  assign n4062 = n2612 & n4034 ;
  assign n4063 = n2613 & n4062 ;
  assign n4064 = ~x114 & n4063 ;
  assign n4065 = n4064 ^ x42 ;
  assign n4103 = n2960 & n4065 ;
  assign n4066 = n4054 ^ n4044 ;
  assign n4067 = n4045 & ~n4047 ;
  assign n4068 = n4066 & n4067 ;
  assign n4069 = n4068 ^ n4045 ;
  assign n4070 = n4069 ^ n2961 ;
  assign n4097 = x219 ^ x199 ;
  assign n4098 = ~n1537 & n4097 ;
  assign n4099 = n4098 ^ x199 ;
  assign n4071 = ~x212 & ~x214 ;
  assign n4072 = n4071 ^ x212 ;
  assign n4073 = n4072 ^ x214 ;
  assign n4083 = x211 & ~x219 ;
  assign n4082 = x219 ^ x211 ;
  assign n4084 = n4083 ^ n4082 ;
  assign n4087 = ~n4073 & ~n4084 ;
  assign n4074 = x199 & ~x200 ;
  assign n4075 = x207 & ~x208 ;
  assign n4076 = n4075 ^ x207 ;
  assign n4077 = ~n4074 & n4076 ;
  assign n4078 = n4077 ^ x200 ;
  assign n4079 = n4078 ^ x211 ;
  assign n4088 = n4087 ^ n4079 ;
  assign n4089 = ~n1537 & n4088 ;
  assign n4090 = n4089 ^ n4078 ;
  assign n4094 = ~n1537 & ~n4083 ;
  assign n4091 = x200 ^ x199 ;
  assign n4092 = n4091 ^ n4074 ;
  assign n4093 = n1537 & ~n4092 ;
  assign n4095 = n4094 ^ n4093 ;
  assign n4096 = ~n4090 & ~n4095 ;
  assign n4100 = n4099 ^ n4096 ;
  assign n4101 = ~n4070 & n4100 ;
  assign n4104 = n4103 ^ n4101 ;
  assign n4112 = ~n4070 & n4090 ;
  assign n4109 = ~x42 & n4064 ;
  assign n4110 = n4109 ^ x43 ;
  assign n4111 = n2960 & n4110 ;
  assign n4114 = n4112 ^ n4111 ;
  assign n4115 = n4052 ^ n4046 ;
  assign n4116 = n4115 ^ x44 ;
  assign n4117 = n4116 ^ n4033 ;
  assign n4118 = n2960 & ~n4117 ;
  assign n4119 = n4115 & ~n4118 ;
  assign n4120 = n4115 ^ n2960 ;
  assign n4121 = n4120 ^ n4118 ;
  assign n4122 = n4121 ^ n4045 ;
  assign n4123 = n4119 & n4122 ;
  assign n4124 = n4123 ^ n4121 ;
  assign n4125 = x979 & n3965 ;
  assign n4127 = n1589 & n1590 ;
  assign n4128 = n1611 & n2759 ;
  assign n4129 = n4127 & n4128 ;
  assign n4130 = ~x24 & n4129 ;
  assign n4131 = n4130 ^ n4129 ;
  assign n4126 = x61 & n3938 ;
  assign n4133 = n4131 ^ n4126 ;
  assign n4144 = n2692 & n3929 ;
  assign n4134 = ~n3936 & ~n3939 ;
  assign n4135 = ~x36 & ~x88 ;
  assign n4136 = ~x104 & ~n2695 ;
  assign n4137 = n4135 & n4136 ;
  assign n4138 = n4137 ^ n2695 ;
  assign n4139 = ~n4134 & ~n4138 ;
  assign n4145 = n4144 ^ n4139 ;
  assign n4146 = ~n3928 & n4145 ;
  assign n4147 = n4146 ^ n4139 ;
  assign n4148 = x48 & n3937 ;
  assign n4185 = n3937 ^ n1337 ;
  assign n4150 = n3937 ^ x49 ;
  assign n4186 = n4185 ^ n4150 ;
  assign n4189 = n4186 ^ x74 ;
  assign n4190 = n4189 ^ n4150 ;
  assign n4187 = n4186 ^ n3248 ;
  assign n4188 = n4187 ^ n4150 ;
  assign n4191 = n4190 ^ n4188 ;
  assign n4168 = ~n3937 & n4150 ;
  assign n4169 = n4189 ^ n4168 ;
  assign n4170 = n4186 ^ n4169 ;
  assign n4171 = n4170 ^ x49 ;
  assign n4195 = n4189 ^ n4188 ;
  assign n4196 = n4195 ^ n4185 ;
  assign n4173 = n4196 ^ x49 ;
  assign n4174 = n4171 & n4173 ;
  assign n4197 = n4196 ^ n3937 ;
  assign n4159 = n4195 ^ n4186 ;
  assign n4175 = n4187 ^ n4159 ;
  assign n4176 = n4197 ^ n4175 ;
  assign n4177 = n4189 ^ n4159 ;
  assign n4178 = n4197 ^ n4177 ;
  assign n4179 = ~n4176 & ~n4178 ;
  assign n4180 = n4174 & n4179 ;
  assign n4181 = n4180 ^ n4168 ;
  assign n4182 = n4191 ^ n4181 ;
  assign n4203 = n4182 ^ n1337 ;
  assign n4204 = n4203 ^ n4197 ;
  assign n4205 = n4204 ^ n4191 ;
  assign n4206 = n4205 ^ n1337 ;
  assign n4207 = n4206 ^ x49 ;
  assign n4208 = n4207 ^ n4197 ;
  assign n4209 = x24 & x50 ;
  assign n4210 = n1745 & n3929 ;
  assign n4211 = ~x86 & n1256 ;
  assign n4212 = ~x58 & n3929 ;
  assign n4213 = n1584 & n4212 ;
  assign n4214 = n4211 & n4213 ;
  assign n4215 = n1245 & n4214 ;
  assign n4216 = ~x94 & x110 ;
  assign n4217 = n4216 ^ n4000 ;
  assign n4218 = n4215 & n4217 ;
  assign n4223 = n3222 ^ n1851 ;
  assign n4226 = x252 & ~n4223 ;
  assign n4227 = n4226 ^ n3222 ;
  assign n4228 = n4218 & ~n4227 ;
  assign n4219 = n3493 ^ n2843 ;
  assign n4220 = n2844 & n3845 ;
  assign n4221 = n4219 & n4220 ;
  assign n4229 = n4228 ^ n4221 ;
  assign n4230 = n4210 & ~n4229 ;
  assign n4231 = n4209 & n4230 ;
  assign n4232 = n4231 ^ n4229 ;
  assign n4233 = n1681 & n1690 ;
  assign n4234 = n1717 & n3935 ;
  assign n4235 = n4233 & n4234 ;
  assign n4236 = n1213 & n4235 ;
  assign n4244 = ~n4070 & ~n4100 ;
  assign n4241 = n2618 & n4033 ;
  assign n4242 = n4241 ^ x52 ;
  assign n4243 = n2960 & n4242 ;
  assign n4248 = n4084 ^ x211 ;
  assign n4249 = ~n4073 & ~n4248 ;
  assign n4250 = n4249 ^ n4082 ;
  assign n4251 = ~n1537 & ~n4250 ;
  assign n4245 = ~x199 & ~n4076 ;
  assign n4246 = n4245 ^ x200 ;
  assign n4247 = n4093 & n4246 ;
  assign n4252 = n4251 ^ n4247 ;
  assign n4253 = ~n4243 & n4252 ;
  assign n4254 = n4244 & n4253 ;
  assign n4255 = n4254 ^ n4243 ;
  assign n4261 = n3965 & n3967 ;
  assign n4256 = n1259 & n2721 ;
  assign n4257 = n4212 & n4256 ;
  assign n4258 = n1594 & n4257 ;
  assign n4259 = ~x24 & n4258 ;
  assign n4260 = n4259 ^ n4258 ;
  assign n4263 = n4261 ^ n4260 ;
  assign n4267 = x106 & n3937 ;
  assign n4266 = x106 & n3936 ;
  assign n4268 = n4267 ^ n4266 ;
  assign n4264 = x24 & n1338 ;
  assign n4265 = n1314 & n4264 ;
  assign n4270 = n4268 ^ n4265 ;
  assign n4272 = x24 & n3835 ;
  assign n4271 = x45 & n3936 ;
  assign n4274 = n4272 ^ n4271 ;
  assign n4275 = x56 ^ x55 ;
  assign n4276 = ~x62 & n4275 ;
  assign n4277 = x841 ^ x24 ;
  assign n4282 = x56 & ~n4277 ;
  assign n4283 = n4282 ^ x24 ;
  assign n4284 = n4276 & ~n4283 ;
  assign n4285 = n1284 & n4284 ;
  assign n4290 = x24 & n1327 ;
  assign n4286 = ~x841 & n1287 ;
  assign n4287 = x62 & x924 ;
  assign n4288 = n4286 & n4287 ;
  assign n4289 = n4288 ^ n4286 ;
  assign n4291 = n4290 ^ n4289 ;
  assign n4292 = n1262 & n2760 ;
  assign n4293 = x841 & n4292 ;
  assign n4294 = n4293 ^ n4292 ;
  assign n4295 = ~x57 & n1289 ;
  assign n4296 = n1283 & n3922 ;
  assign n4297 = n4295 & n4296 ;
  assign n4298 = n4297 ^ n4288 ;
  assign n4299 = n3965 & n3969 ;
  assign n4300 = n1246 & n4257 ;
  assign n4301 = ~x24 & n4300 ;
  assign n4302 = n4301 ^ n4300 ;
  assign n4303 = ~n4299 & ~n4302 ;
  assign n4304 = x61 & n3937 ;
  assign n4305 = n4304 ^ n4301 ;
  assign n4306 = x62 ^ x57 ;
  assign n4307 = ~n1341 & n4306 ;
  assign n4310 = x62 & ~n4277 ;
  assign n4311 = n4310 ^ x24 ;
  assign n4312 = n4307 & ~n4311 ;
  assign n4313 = x63 & n3939 ;
  assign n4314 = ~x999 & n4313 ;
  assign n4315 = n4314 ^ n4313 ;
  assign n4316 = ~n4130 & ~n4315 ;
  assign n4317 = x107 & n3939 ;
  assign n4319 = n4317 ^ n3941 ;
  assign n4320 = n3965 & n3974 ;
  assign n4321 = ~n3972 & n4320 ;
  assign n4322 = x299 & n4097 ;
  assign n4323 = n4322 ^ x199 ;
  assign n4324 = x81 & x314 ;
  assign n4325 = n1621 & n3935 ;
  assign n4326 = n1243 & n4325 ;
  assign n4327 = n4324 & n4326 ;
  assign n4328 = n4323 & n4327 ;
  assign n4329 = ~x69 & n1709 ;
  assign n4330 = n4234 & n4329 ;
  assign n4331 = x314 & n4330 ;
  assign n4332 = x83 & ~x103 ;
  assign n4333 = n4331 & n4332 ;
  assign n4334 = n2824 & n2966 ;
  assign n4337 = n1936 & ~n2672 ;
  assign n4335 = x299 & n1350 ;
  assign n4336 = ~n2686 & n4335 ;
  assign n4338 = n4337 ^ n4336 ;
  assign n4339 = n4334 & n4338 ;
  assign n4340 = ~x71 & n3936 ;
  assign n4341 = ~x314 & n4340 ;
  assign n4342 = x69 & n4341 ;
  assign n4343 = n4342 ^ n4340 ;
  assign n4344 = n4343 ^ n3936 ;
  assign n4345 = n2654 & n2966 ;
  assign n4346 = ~n4334 & ~n4345 ;
  assign n4349 = n1424 & ~n2672 ;
  assign n4350 = x198 & n4349 ;
  assign n4347 = n1511 & ~n2686 ;
  assign n4348 = x210 & n4347 ;
  assign n4351 = n4350 ^ n4348 ;
  assign n4352 = x589 & n4351 ;
  assign n4353 = ~n4346 & n4352 ;
  assign n4354 = x593 & n4353 ;
  assign n4355 = n4354 ^ n4353 ;
  assign n4356 = ~x24 & x70 ;
  assign n4357 = n4356 ^ x70 ;
  assign n4359 = n2792 & n4357 ;
  assign n4360 = n4359 ^ n3964 ;
  assign n4361 = ~n4355 & ~n4360 ;
  assign n4362 = n4092 ^ x199 ;
  assign n4363 = n4362 ^ n4248 ;
  assign n4364 = ~x299 & n4363 ;
  assign n4365 = n4364 ^ n4248 ;
  assign n4366 = n4365 ^ n4323 ;
  assign n4375 = n4327 & n4366 ;
  assign n4367 = ~n1706 & n4234 ;
  assign n4368 = x85 & ~n1232 ;
  assign n4369 = n1662 & n1667 ;
  assign n4370 = n4368 & n4369 ;
  assign n4371 = ~x314 & n4370 ;
  assign n4372 = n4371 ^ n4370 ;
  assign n4373 = n4367 & n4372 ;
  assign n4376 = n4375 ^ n4373 ;
  assign n4377 = n3238 & n4334 ;
  assign n4378 = ~x38 & x88 ;
  assign n4379 = n1762 & n2696 ;
  assign n4380 = n4378 & n4379 ;
  assign n4381 = n4380 ^ x38 ;
  assign n4382 = n1556 & ~n4381 ;
  assign n4386 = x72 & n1757 ;
  assign n4391 = n4382 & n4386 ;
  assign n4392 = x24 & n4391 ;
  assign n4393 = n4392 ^ x24 ;
  assign n4383 = n4382 ^ n1556 ;
  assign n4384 = n4383 ^ x24 ;
  assign n4394 = n4393 ^ n4384 ;
  assign n4395 = ~n4377 & ~n4394 ;
  assign n4396 = x314 & x1050 ;
  assign n4397 = n4396 ^ x1050 ;
  assign n4398 = ~x39 & ~n4397 ;
  assign n4400 = n2688 & n4334 ;
  assign n4399 = x73 & n1919 ;
  assign n4402 = n4400 ^ n4399 ;
  assign n4403 = n4398 & n4402 ;
  assign n4404 = n4403 ^ n4402 ;
  assign n4417 = x74 & n4264 ;
  assign n4405 = n1556 & ~n1851 ;
  assign n4409 = ~x479 & ~x841 ;
  assign n4406 = x479 & n1784 ;
  assign n4407 = n2608 & n4406 ;
  assign n4408 = n4407 ^ n2608 ;
  assign n4410 = n4409 ^ n4408 ;
  assign n4413 = ~x96 & n4410 ;
  assign n4414 = n4413 ^ n4409 ;
  assign n4415 = n4405 & n4414 ;
  assign n4416 = n1860 & n4415 ;
  assign n4419 = n4417 ^ n4416 ;
  assign n4421 = x75 & n4264 ;
  assign n4420 = n1556 & n1871 ;
  assign n4423 = n4421 ^ n4420 ;
  assign n4424 = n3455 & ~n3889 ;
  assign n4431 = n3198 & n3459 ;
  assign n4425 = n3222 ^ x94 ;
  assign n4426 = n4425 ^ n4424 ;
  assign n4432 = n4431 ^ n4426 ;
  assign n4433 = n4424 & n4432 ;
  assign n4434 = n4433 ^ n4426 ;
  assign n4435 = n4434 ^ x94 ;
  assign n4436 = n4434 ^ n3222 ;
  assign n4437 = ~n4433 & ~n4436 ;
  assign n4438 = ~n4435 & n4437 ;
  assign n4439 = n4438 ^ n4434 ;
  assign n4440 = n1851 & ~n4439 ;
  assign n4441 = n3459 ^ x252 ;
  assign n4444 = x94 & n4441 ;
  assign n4445 = n4444 ^ n3459 ;
  assign n4446 = n4440 & n4445 ;
  assign n4447 = n4446 ^ n4439 ;
  assign n4448 = n1919 & ~n4447 ;
  assign n4449 = x77 & x314 ;
  assign n4450 = n4449 ^ n1257 ;
  assign n4451 = n2792 & ~n4450 ;
  assign n4452 = x232 & n3000 ;
  assign n4468 = x182 ^ x160 ;
  assign n4469 = ~x299 & n4468 ;
  assign n4470 = n4469 ^ x160 ;
  assign n4471 = n2806 & n3219 ;
  assign n4472 = ~n4470 & n4471 ;
  assign n4479 = n4472 ^ n3620 ;
  assign n4453 = ~x166 & n3539 ;
  assign n4454 = n3618 & n4453 ;
  assign n4455 = n4454 ^ x163 ;
  assign n4456 = ~x163 & ~n4455 ;
  assign n4457 = x299 & n4456 ;
  assign n4458 = ~n3631 & ~n4457 ;
  assign n4459 = x153 & n1607 ;
  assign n4460 = n2811 & n4459 ;
  assign n4461 = n4460 ^ n1765 ;
  assign n4462 = ~n1765 & ~n4461 ;
  assign n4463 = n1810 & ~n4462 ;
  assign n4464 = n4463 ^ x175 ;
  assign n4465 = x299 & n4464 ;
  assign n4466 = n4465 ^ x175 ;
  assign n4467 = ~n4458 & ~n4466 ;
  assign n4473 = n4472 ^ n3219 ;
  assign n4474 = ~n4467 & n4473 ;
  assign n4480 = x189 ^ x166 ;
  assign n4481 = ~x299 & n4480 ;
  assign n4482 = n4481 ^ x166 ;
  assign n4483 = n4474 & n4482 ;
  assign n4484 = n4479 & n4483 ;
  assign n4475 = ~x34 & n3713 ;
  assign n4476 = n4475 ^ x79 ;
  assign n4477 = n4476 ^ n3549 ;
  assign n4478 = n4477 ^ n4474 ;
  assign n4485 = n4484 ^ n4478 ;
  assign n4486 = n4485 ^ n4477 ;
  assign n4494 = ~x184 & n4486 ;
  assign n4495 = ~n3673 & n4494 ;
  assign n4496 = n4495 ^ n3673 ;
  assign n4488 = n4485 ^ n3673 ;
  assign n4497 = n4496 ^ n4488 ;
  assign n4498 = ~n3626 & ~n4497 ;
  assign n4499 = n4498 ^ n4477 ;
  assign n4500 = ~x39 & n4499 ;
  assign n4501 = ~x38 & n3210 ;
  assign n4503 = ~x166 & n3585 ;
  assign n4502 = ~x189 & n3583 ;
  assign n4504 = n4503 ^ n4502 ;
  assign n4505 = n2824 & n4504 ;
  assign n4507 = x156 & n3585 ;
  assign n4506 = x179 & n3583 ;
  assign n4508 = n4507 ^ n4506 ;
  assign n4509 = n2654 & n4508 ;
  assign n4510 = ~n4505 & ~n4509 ;
  assign n4511 = n3219 & ~n4510 ;
  assign n4512 = n3537 & n4511 ;
  assign n4513 = x39 & ~n4512 ;
  assign n4514 = n3539 & n4513 ;
  assign n4517 = n4514 ^ n3539 ;
  assign n4515 = ~n3602 & ~n4477 ;
  assign n4516 = n4514 & n4515 ;
  assign n4518 = n4517 ^ n4516 ;
  assign n4519 = n4501 & n4518 ;
  assign n4520 = ~n4500 & n4519 ;
  assign n4521 = n1450 & n3539 ;
  assign n4522 = x179 ^ x156 ;
  assign n4525 = x299 & n4522 ;
  assign n4526 = n4525 ^ x179 ;
  assign n4527 = n3219 & n4526 ;
  assign n4528 = n4527 ^ n4477 ;
  assign n4531 = n3735 & ~n4528 ;
  assign n4532 = n4531 ^ n4477 ;
  assign n4533 = n4521 & ~n4532 ;
  assign n4534 = n4533 ^ n1450 ;
  assign n4535 = ~n1307 & ~n4534 ;
  assign n4536 = ~x40 & ~n3575 ;
  assign n4537 = ~n4535 & n4536 ;
  assign n4538 = ~n4520 & n4537 ;
  assign n4539 = n1449 & n3219 ;
  assign n4540 = x187 ^ x147 ;
  assign n4543 = ~x299 & n4540 ;
  assign n4544 = n4543 ^ x147 ;
  assign n4545 = n4539 & n4544 ;
  assign n4546 = n4545 ^ n1449 ;
  assign n4547 = n1275 & n3219 ;
  assign n4552 = n3786 ^ x145 ;
  assign n4553 = n3788 & n4552 ;
  assign n4554 = n4553 ^ x140 ;
  assign n4555 = n4554 ^ x184 ;
  assign n4548 = n3783 ^ x197 ;
  assign n4549 = n3784 & n4548 ;
  assign n4550 = n4549 ^ x162 ;
  assign n4551 = n4550 ^ x163 ;
  assign n4556 = n4555 ^ n4551 ;
  assign n4559 = ~x299 & n4556 ;
  assign n4560 = n4559 ^ n4551 ;
  assign n4561 = n4547 & n4560 ;
  assign n4562 = ~n4546 & ~n4561 ;
  assign n4563 = ~n4538 & n4562 ;
  assign n4564 = n1290 & ~n4563 ;
  assign n4565 = ~n1290 & ~n3702 ;
  assign n4570 = ~x147 & ~n1275 ;
  assign n4566 = n3219 ^ n1275 ;
  assign n4571 = n4570 ^ n4566 ;
  assign n4572 = n4551 ^ x74 ;
  assign n4573 = ~n1275 & ~n4572 ;
  assign n4574 = n4573 ^ n4551 ;
  assign n4575 = n4566 & n4574 ;
  assign n4576 = n4571 & n4575 ;
  assign n4577 = n4576 ^ n4573 ;
  assign n4578 = n4577 ^ n4551 ;
  assign n4579 = n4565 & n4578 ;
  assign n4580 = ~x40 & ~n1289 ;
  assign n4583 = x163 & n3219 ;
  assign n4584 = n4583 ^ n4477 ;
  assign n4585 = n3718 & ~n4584 ;
  assign n4586 = n4585 ^ n4477 ;
  assign n4587 = n3539 & ~n4586 ;
  assign n4588 = n3702 & ~n4587 ;
  assign n4589 = n4580 & n4588 ;
  assign n4590 = ~n4579 & ~n4589 ;
  assign n4591 = ~n4564 & n4590 ;
  assign n4601 = x98 & ~x592 ;
  assign n4602 = x1199 & n4601 ;
  assign n4595 = ~x592 & ~n3034 ;
  assign n4596 = n3188 & n4595 ;
  assign n4597 = n4596 ^ n3188 ;
  assign n4592 = ~x588 & ~x590 ;
  assign n4593 = n4592 ^ n3351 ;
  assign n4594 = n4593 ^ n2958 ;
  assign n4598 = n3200 ^ x590 ;
  assign n4599 = ~n3198 & ~n4598 ;
  assign n4600 = n4599 ^ x590 ;
  assign n4603 = n4602 ^ n3198 ;
  assign n4604 = n4603 ^ n4597 ;
  assign n4605 = ~n4600 & ~n4604 ;
  assign n4606 = n4605 ^ n3198 ;
  assign n4607 = n4597 & ~n4606 ;
  assign n4608 = n4607 ^ n4592 ;
  assign n4609 = n4608 ^ n2958 ;
  assign n4610 = n4607 ^ n3186 ;
  assign n4611 = n4610 ^ n3351 ;
  assign n4612 = ~n4609 & n4611 ;
  assign n4613 = ~n4594 & n4612 ;
  assign n4614 = n4613 ^ n4607 ;
  assign n4615 = n4614 ^ n3351 ;
  assign n4616 = n2958 & n4615 ;
  assign n4617 = n3351 & n4616 ;
  assign n4618 = n3320 & n4617 ;
  assign n4619 = ~x63 & n1341 ;
  assign n4620 = ~n2761 & n4619 ;
  assign n4621 = n4620 ^ n1341 ;
  assign n4622 = n4618 & ~n4621 ;
  assign n4623 = n3201 & ~n4622 ;
  assign n4631 = n4597 & n4623 ;
  assign n4632 = ~n4602 & n4631 ;
  assign n4633 = n4632 ^ n4602 ;
  assign n4624 = n4623 ^ n4622 ;
  assign n4625 = n4624 ^ n4602 ;
  assign n4634 = n4633 ^ n4625 ;
  assign n4635 = n3167 & n4634 ;
  assign n4636 = ~n3207 & ~n4635 ;
  assign n4637 = ~x80 & n3209 ;
  assign n4638 = ~n4636 & n4637 ;
  assign n4639 = ~x68 & ~n4134 ;
  assign n4640 = ~x314 & n4639 ;
  assign n4641 = x81 & n4640 ;
  assign n4642 = n4641 ^ n4639 ;
  assign n4643 = n4642 ^ n4134 ;
  assign n4644 = x314 ^ x66 ;
  assign n4647 = ~x69 & n4644 ;
  assign n4648 = n4647 ^ x314 ;
  assign n4649 = n3936 & n4648 ;
  assign n4653 = ~x314 & n4330 ;
  assign n4654 = n4332 & n4653 ;
  assign n4650 = ~x68 & x84 ;
  assign n4651 = n1244 & n4367 ;
  assign n4652 = n4650 & n4651 ;
  assign n4655 = n4654 ^ n4652 ;
  assign n4656 = n4327 & ~n4365 ;
  assign n4657 = ~x67 & n4367 ;
  assign n4658 = ~n4371 & n4657 ;
  assign n4659 = n4658 ^ n4367 ;
  assign n4660 = n4338 & n4345 ;
  assign n4661 = n2781 & n4331 ;
  assign n4662 = x88 & n2607 ;
  assign n4668 = n3939 & n4662 ;
  assign n4663 = x104 & n2695 ;
  assign n4664 = n3936 & n4663 ;
  assign n4665 = ~n3198 & n4664 ;
  assign n4666 = n4665 ^ n4664 ;
  assign n4669 = n4668 ^ n4666 ;
  assign n4670 = n2792 & ~n4356 ;
  assign n4671 = x89 & n4670 ;
  assign n4672 = x841 & n4671 ;
  assign n4673 = n4672 ^ n4670 ;
  assign n4674 = n4673 ^ n2792 ;
  assign n4675 = ~x1050 & n4399 ;
  assign n4676 = n4675 ^ n4293 ;
  assign n4685 = n2966 & n3239 ;
  assign n4677 = n3292 ^ n1864 ;
  assign n4678 = n4677 ^ n4212 ;
  assign n4679 = n3927 ^ x24 ;
  assign n4680 = n1864 & ~n4679 ;
  assign n4681 = n4680 ^ x24 ;
  assign n4682 = ~n4678 & n4681 ;
  assign n4683 = n4682 ^ n1864 ;
  assign n4684 = n4212 & n4683 ;
  assign n4687 = n4685 ^ n4684 ;
  assign n4690 = x92 & n4397 ;
  assign n4691 = n4690 ^ n2689 ;
  assign n4692 = ~x39 & n4691 ;
  assign n4693 = n4692 ^ n2689 ;
  assign n4694 = n1303 & n4693 ;
  assign n4696 = n1328 & n1451 ;
  assign n4697 = ~x1050 & n4696 ;
  assign n4695 = n2717 & n2792 ;
  assign n4699 = n4697 ^ n4695 ;
  assign n4736 = n3938 ^ n3250 ;
  assign n4701 = n3938 ^ x49 ;
  assign n4737 = n4736 ^ n4701 ;
  assign n4740 = n4737 ^ n4218 ;
  assign n4741 = n4740 ^ n4701 ;
  assign n4738 = n4737 ^ n1851 ;
  assign n4739 = n4738 ^ n4701 ;
  assign n4742 = n4741 ^ n4739 ;
  assign n4746 = n4740 ^ n4739 ;
  assign n4747 = n4746 ^ n4736 ;
  assign n4748 = n4747 ^ n3938 ;
  assign n4719 = ~n3938 & n4701 ;
  assign n4720 = n4740 ^ n4719 ;
  assign n4721 = n4737 ^ n4720 ;
  assign n4722 = n4721 ^ x49 ;
  assign n4724 = n4747 ^ x49 ;
  assign n4725 = n4722 & ~n4724 ;
  assign n4710 = n4746 ^ n4737 ;
  assign n4726 = n4738 ^ n4710 ;
  assign n4727 = n4748 ^ n4726 ;
  assign n4728 = n4740 ^ n4710 ;
  assign n4729 = n4748 ^ n4728 ;
  assign n4730 = n4727 & ~n4729 ;
  assign n4731 = n4725 & n4730 ;
  assign n4732 = n4731 ^ n4719 ;
  assign n4733 = n4742 ^ n4732 ;
  assign n4734 = n4733 ^ n3250 ;
  assign n4735 = n4748 ^ n4734 ;
  assign n4743 = n4742 ^ n4735 ;
  assign n4751 = n4743 ^ n3250 ;
  assign n4752 = n4751 ^ x49 ;
  assign n4753 = n4752 ^ n4748 ;
  assign n4816 = ~x32 & ~x40 ;
  assign n4817 = n1556 & n4816 ;
  assign n4818 = x95 & n1270 ;
  assign n4819 = n4817 & n4818 ;
  assign n4820 = x24 & n4819 ;
  assign n4755 = n4349 ^ n4347 ;
  assign n4756 = ~n4346 & n4755 ;
  assign n4792 = n4756 ^ n3938 ;
  assign n4757 = n4756 ^ n4352 ;
  assign n4793 = n4792 ^ n4757 ;
  assign n4796 = n4793 ^ x89 ;
  assign n4797 = n4796 ^ n4757 ;
  assign n4794 = n4793 ^ x332 ;
  assign n4795 = n4794 ^ n4757 ;
  assign n4798 = n4797 ^ n4795 ;
  assign n4775 = ~n4756 & ~n4757 ;
  assign n4776 = n4794 ^ n4775 ;
  assign n4777 = n4793 ^ n4776 ;
  assign n4778 = n4777 ^ n4352 ;
  assign n4802 = n4796 ^ n4795 ;
  assign n4803 = n4802 ^ n4792 ;
  assign n4780 = n4803 ^ n4352 ;
  assign n4781 = n4778 & ~n4780 ;
  assign n4804 = n4803 ^ n4756 ;
  assign n4766 = n4802 ^ n4793 ;
  assign n4782 = n4796 ^ n4766 ;
  assign n4783 = n4804 ^ n4782 ;
  assign n4784 = n4794 ^ n4766 ;
  assign n4785 = n4804 ^ n4784 ;
  assign n4786 = ~n4783 & n4785 ;
  assign n4787 = n4781 & n4786 ;
  assign n4788 = n4787 ^ n4775 ;
  assign n4789 = n4798 ^ n4788 ;
  assign n4810 = n4789 ^ n3938 ;
  assign n4811 = n4810 ^ n4804 ;
  assign n4812 = n4811 ^ n4798 ;
  assign n4813 = n4812 ^ n3938 ;
  assign n4814 = n4813 ^ n4352 ;
  assign n4815 = n4814 ^ n4804 ;
  assign n4822 = n4820 ^ n4815 ;
  assign n4823 = x96 ^ x95 ;
  assign n4826 = ~n1852 & ~n4409 ;
  assign n4827 = n4826 ^ x24 ;
  assign n4828 = x96 & ~n4827 ;
  assign n4829 = n4828 ^ x24 ;
  assign n4830 = n4823 & ~n4829 ;
  assign n4831 = n4817 & n4830 ;
  assign n4832 = ~n1270 & n4831 ;
  assign n4833 = ~n1762 & n4832 ;
  assign n4834 = n4833 ^ n4831 ;
  assign n4835 = n1857 & ~n1864 ;
  assign n4836 = n3929 & ~n4408 ;
  assign n4837 = n4835 & n4836 ;
  assign n4838 = ~n4354 & ~n4837 ;
  assign n4839 = n4696 ^ n4399 ;
  assign n4840 = n4396 & n4839 ;
  assign n4850 = n4056 ^ n4049 ;
  assign n4849 = ~x144 & n4056 ;
  assign n4851 = n4850 ^ n4849 ;
  assign n4848 = ~x161 & n4049 ;
  assign n4852 = n4851 ^ n4848 ;
  assign n4853 = n4045 & n4852 ;
  assign n4845 = n2610 & n4034 ;
  assign n4846 = n4845 ^ x99 ;
  assign n4847 = n2960 & n4846 ;
  assign n4854 = n4853 ^ n4847 ;
  assign n4855 = x683 ^ x252 ;
  assign n4856 = ~n1797 & ~n4855 ;
  assign n4857 = n4856 ^ x683 ;
  assign n4858 = ~n3222 & n3485 ;
  assign n4859 = ~n4857 & n4858 ;
  assign n4867 = n4856 & n4859 ;
  assign n4868 = n2695 & n4867 ;
  assign n4869 = n4868 ^ n2695 ;
  assign n4860 = n4859 ^ n3485 ;
  assign n4861 = n4860 ^ n2695 ;
  assign n4870 = n4869 ^ n4861 ;
  assign n4871 = n1274 & ~n4870 ;
  assign n4872 = n2844 & ~n4871 ;
  assign n4874 = ~n3249 & n3492 ;
  assign n4875 = n4872 & n4874 ;
  assign n4873 = n4872 ^ n2844 ;
  assign n4876 = n4875 ^ n4873 ;
  assign n4877 = n4849 ^ n4848 ;
  assign n4881 = n4045 & n4877 ;
  assign n4878 = n4034 ^ x101 ;
  assign n4879 = n2960 & n4878 ;
  assign n4882 = n4881 ^ n4879 ;
  assign n4883 = x65 & n3939 ;
  assign n4885 = n4215 & n4216 ;
  assign n4886 = n2695 & ~n3222 ;
  assign n4887 = n4885 & n4886 ;
  assign n4888 = n4887 ^ n4885 ;
  assign n4889 = ~n4665 & ~n4888 ;
  assign n4890 = n4267 ^ n4259 ;
  assign n4892 = n3953 ^ x108 ;
  assign n4893 = ~x98 & n4210 ;
  assign n4894 = ~n4892 & n4893 ;
  assign n4895 = n4894 ^ n4210 ;
  assign n4891 = n2964 & ~n4621 ;
  assign n4897 = n4895 ^ n4891 ;
  assign n4898 = n4210 & n4449 ;
  assign n4899 = n2781 & n4235 ;
  assign n4900 = ~x314 & n4899 ;
  assign n4901 = n4900 ^ n4899 ;
  assign n4902 = ~n4887 & ~n4901 ;
  assign n4903 = ~x24 & n1556 ;
  assign n4905 = n4386 & n4903 ;
  assign n4906 = n4905 ^ n4900 ;
  assign n4907 = x124 & ~x468 ;
  assign n4912 = n2611 & n4034 ;
  assign n4913 = n4912 ^ x113 ;
  assign n4914 = n2960 & n4913 ;
  assign n4915 = n4063 ^ x114 ;
  assign n4916 = n2960 & n4915 ;
  assign n4921 = ~x116 & n4062 ;
  assign n4922 = n4921 ^ x115 ;
  assign n4923 = n2960 & n4922 ;
  assign n4924 = n4062 ^ x116 ;
  assign n4925 = n2960 & n4924 ;
  assign n4926 = x87 & n3219 ;
  assign n4927 = n4926 ^ n3219 ;
  assign n4928 = n3537 & n4927 ;
  assign n4933 = x178 & n2654 ;
  assign n4932 = x190 & n2824 ;
  assign n4934 = n4933 ^ n4932 ;
  assign n4935 = n3583 & n4934 ;
  assign n4937 = x157 & n2654 ;
  assign n4936 = x168 & n2824 ;
  assign n4938 = n4937 ^ n4936 ;
  assign n4939 = n3585 & n4938 ;
  assign n4940 = ~n4935 & ~n4939 ;
  assign n4929 = x178 ^ x157 ;
  assign n4930 = ~x299 & n4929 ;
  assign n4931 = n4930 ^ x157 ;
  assign n4941 = n4940 ^ n4931 ;
  assign n4944 = x92 & ~n4941 ;
  assign n4945 = n4944 ^ n4940 ;
  assign n4946 = n1298 & ~n4945 ;
  assign n4947 = n4928 & n4946 ;
  assign n4948 = n3540 & ~n4947 ;
  assign n4976 = n1282 & ~n3626 ;
  assign n4977 = n3219 & n3631 ;
  assign n4978 = x173 ^ x151 ;
  assign n4981 = ~x299 & n4978 ;
  assign n4982 = n4981 ^ x151 ;
  assign n4983 = n4977 & ~n4982 ;
  assign n4984 = n4983 ^ n3219 ;
  assign n4985 = ~n2806 & ~n4984 ;
  assign n4986 = ~x150 & x299 ;
  assign n4987 = ~n3645 & n4986 ;
  assign n4988 = n4987 ^ x299 ;
  assign n4990 = x73 & ~x168 ;
  assign n4991 = n4988 & n4990 ;
  assign n4992 = n4991 ^ n4987 ;
  assign n4993 = ~x185 & ~x299 ;
  assign n4994 = ~x73 & x232 ;
  assign n4995 = ~n1780 & n3645 ;
  assign n4996 = n4994 & n4995 ;
  assign n4997 = n4996 ^ n3645 ;
  assign n4998 = n4993 & ~n4997 ;
  assign n4999 = n4998 ^ x299 ;
  assign n5002 = n4998 ^ x190 ;
  assign n5003 = x73 & ~n5002 ;
  assign n5004 = ~n4999 & n5003 ;
  assign n5005 = n5004 ^ n4999 ;
  assign n5006 = n5005 ^ x299 ;
  assign n5007 = ~n4992 & ~n5006 ;
  assign n5008 = ~n4985 & n5007 ;
  assign n4949 = ~x54 & n1448 ;
  assign n4950 = x39 ^ x38 ;
  assign n4951 = ~x92 & n4950 ;
  assign n4952 = ~x38 & n4951 ;
  assign n4953 = ~n3601 & n4952 ;
  assign n4954 = n4953 ^ n4951 ;
  assign n4955 = n4954 ^ x92 ;
  assign n4956 = n4949 & n4955 ;
  assign n4957 = n1273 & n4956 ;
  assign n4967 = ~n1311 & ~n3210 ;
  assign n4961 = n4957 ^ n1450 ;
  assign n4959 = n3549 ^ x118 ;
  assign n4958 = ~x79 & n4475 ;
  assign n4960 = n4959 ^ n4958 ;
  assign n4962 = n4961 ^ n4960 ;
  assign n4968 = n4967 ^ n4962 ;
  assign n4969 = n4957 & n4968 ;
  assign n4970 = n4969 ^ n4962 ;
  assign n4971 = n4970 ^ n1450 ;
  assign n4972 = n4970 ^ n4957 ;
  assign n4973 = ~n4969 & ~n4972 ;
  assign n4974 = ~n4971 & n4973 ;
  assign n4975 = n4974 ^ n4970 ;
  assign n5009 = n5008 ^ n4975 ;
  assign n5010 = n4976 & n5009 ;
  assign n5011 = n5010 ^ n4975 ;
  assign n5012 = n4948 & ~n5011 ;
  assign n5013 = n3219 ^ n1289 ;
  assign n5014 = n1289 & ~n1537 ;
  assign n5023 = x165 & n3701 ;
  assign n5024 = n3219 & n5023 ;
  assign n5025 = n5024 ^ n3701 ;
  assign n5019 = ~x163 & ~n4550 ;
  assign n5020 = n5019 ^ x150 ;
  assign n5021 = n4547 & ~n5020 ;
  assign n5026 = n5025 ^ n5021 ;
  assign n5027 = n5014 & n5026 ;
  assign n5028 = n5027 ^ n1289 ;
  assign n5029 = n3701 & n5028 ;
  assign n5030 = n5013 & n5029 ;
  assign n5031 = n5030 ^ n5028 ;
  assign n5032 = ~x299 & n4547 ;
  assign n5037 = ~x184 & ~n4554 ;
  assign n5038 = n5037 ^ x185 ;
  assign n5039 = n5032 & ~n5038 ;
  assign n5040 = n5039 ^ x299 ;
  assign n5048 = ~x143 & ~n5040 ;
  assign n5049 = n1449 & n5048 ;
  assign n5050 = n5049 ^ n1449 ;
  assign n5042 = n5039 ^ n1449 ;
  assign n5051 = n5050 ^ n5042 ;
  assign n5052 = n5031 & ~n5051 ;
  assign n5053 = ~n5012 & n5052 ;
  assign n5056 = x150 & n3219 ;
  assign n5057 = n5056 ^ n4960 ;
  assign n5058 = n1325 & ~n5057 ;
  assign n5059 = n5058 ^ n4960 ;
  assign n5060 = n3703 & ~n5059 ;
  assign n5061 = n5060 ^ n3703 ;
  assign n5062 = ~n1290 & ~n5061 ;
  assign n5063 = ~n5026 & n5062 ;
  assign n5064 = ~n5053 & ~n5063 ;
  assign n5082 = n3237 & n4345 ;
  assign n5065 = n1465 & n2844 ;
  assign n5066 = n1866 ^ n1257 ;
  assign n5067 = n5066 ^ n1607 ;
  assign n5068 = n1605 & ~n2758 ;
  assign n5069 = n5068 ^ n1257 ;
  assign n5070 = n5069 ^ n1607 ;
  assign n5071 = n5068 ^ x109 ;
  assign n5072 = n5071 ^ n1866 ;
  assign n5073 = n5070 & n5072 ;
  assign n5074 = ~n5067 & n5073 ;
  assign n5075 = n5074 ^ n5068 ;
  assign n5076 = n5075 ^ n1866 ;
  assign n5077 = n1607 & ~n5076 ;
  assign n5078 = ~n1866 & n5077 ;
  assign n5079 = n1919 & ~n5078 ;
  assign n5080 = ~n4696 & ~n5079 ;
  assign n5081 = ~n5065 & n5080 ;
  assign n5084 = n5082 ^ n5081 ;
  assign n5085 = n5084 ^ x128 ;
  assign n5086 = ~x228 & ~n5085 ;
  assign n5087 = n5086 ^ x128 ;
  assign n5088 = ~x31 & ~x80 ;
  assign n5089 = x818 & n5088 ;
  assign n5090 = x951 & x982 ;
  assign n5091 = n3009 & n3209 ;
  assign n5092 = n5090 & n5091 ;
  assign n5093 = ~n5089 & ~n5092 ;
  assign n5094 = n1290 & ~n3201 ;
  assign n5095 = ~n3333 & n5094 ;
  assign n5096 = n5095 ^ n3201 ;
  assign n5097 = ~x120 & ~n5096 ;
  assign n5098 = ~n5093 & n5097 ;
  assign n5099 = x1093 & n5098 ;
  assign n5100 = n5099 ^ n5097 ;
  assign n5101 = n5100 ^ n5096 ;
  assign n5102 = n2832 & n3810 ;
  assign n5123 = n3965 & n5102 ;
  assign n5108 = x184 ^ x163 ;
  assign n5109 = n1537 & n5108 ;
  assign n5110 = n5109 ^ x163 ;
  assign n5105 = ~n1537 & n1794 ;
  assign n5106 = n5105 ^ x142 ;
  assign n5107 = x51 & n5106 ;
  assign n5111 = n5110 ^ n5107 ;
  assign n5112 = ~x87 & ~n5111 ;
  assign n5113 = n5112 ^ n5110 ;
  assign n5114 = ~n1209 & ~n2964 ;
  assign n5117 = n1537 & n3796 ;
  assign n5118 = n5117 ^ x161 ;
  assign n5119 = n5114 & n5118 ;
  assign n5120 = n5119 ^ n2965 ;
  assign n5121 = n5113 & ~n5120 ;
  assign n5124 = n5123 ^ n5121 ;
  assign n5125 = ~x24 & n4449 ;
  assign n5126 = n2792 & n3658 ;
  assign n5127 = n5125 & n5126 ;
  assign n5128 = n5127 ^ n3219 ;
  assign n5129 = n3219 & n5128 ;
  assign n5130 = ~n5124 & n5129 ;
  assign n5131 = n5130 ^ n3219 ;
  assign n5132 = ~x39 & n1855 ;
  assign n5133 = ~x24 & x77 ;
  assign n5134 = n5133 ^ x77 ;
  assign n5135 = ~x86 & ~n5134 ;
  assign n5136 = ~n4449 & n5135 ;
  assign n5137 = n2958 & ~n5136 ;
  assign n5138 = n5132 & n5137 ;
  assign n5139 = n1736 & n5138 ;
  assign n5159 = n4527 & ~n5125 ;
  assign n5140 = x72 ^ x39 ;
  assign n5141 = n2959 & n5140 ;
  assign n5142 = x39 & ~n2825 ;
  assign n5143 = n5141 & n5142 ;
  assign n5144 = n5143 ^ n5141 ;
  assign n5147 = ~x134 & ~x135 ;
  assign n5148 = ~x136 & n5147 ;
  assign n5145 = ~x125 & ~x133 ;
  assign n5149 = ~x121 & n5145 ;
  assign n5150 = x126 & ~x132 ;
  assign n5151 = n5150 ^ x132 ;
  assign n5152 = n5149 & ~n5151 ;
  assign n5153 = ~x130 & n5152 ;
  assign n5154 = n5148 & n5153 ;
  assign n5146 = n5145 ^ x121 ;
  assign n5155 = n5154 ^ n5146 ;
  assign n5156 = ~n5144 & ~n5155 ;
  assign n5160 = n5159 ^ n5156 ;
  assign n5161 = n5139 & n5160 ;
  assign n5162 = n5161 ^ n5156 ;
  assign n5163 = n2965 & n5162 ;
  assign n5164 = ~n5131 & ~n5163 ;
  assign n5165 = ~x72 & ~x90 ;
  assign n5166 = ~x111 & n2779 ;
  assign n5167 = n5165 & n5166 ;
  assign n5168 = n2792 & ~n5167 ;
  assign n5170 = ~x39 & x110 ;
  assign n5173 = ~n2619 & n2695 ;
  assign n5174 = n5170 & n5173 ;
  assign n5183 = n4115 & n5174 ;
  assign n5184 = n3219 & n5183 ;
  assign n5185 = n5184 ^ n3219 ;
  assign n5169 = x110 ^ x39 ;
  assign n5171 = n5170 ^ n5169 ;
  assign n5172 = n2976 & n5171 ;
  assign n5175 = n5174 ^ n5172 ;
  assign n5176 = n5175 ^ n3219 ;
  assign n5186 = n5185 ^ n5176 ;
  assign n5187 = ~n5168 & ~n5186 ;
  assign n5196 = ~x152 & ~n1209 ;
  assign n5197 = n5196 ^ x172 ;
  assign n5198 = ~x51 & n5197 ;
  assign n5199 = n5198 ^ x172 ;
  assign n5226 = x299 & n3219 ;
  assign n5227 = ~n5199 & n5226 ;
  assign n5228 = n5227 ^ n3219 ;
  assign n5243 = ~x287 & n3219 ;
  assign n5244 = x158 & n1347 ;
  assign n5245 = n5243 & n5244 ;
  assign n5246 = n5245 ^ n1273 ;
  assign n5247 = n1273 & n5246 ;
  assign n5248 = ~n3233 & n5247 ;
  assign n5249 = n5248 ^ n1273 ;
  assign n5250 = ~n5228 & ~n5249 ;
  assign n5231 = ~x174 & ~n1209 ;
  assign n5232 = n5231 ^ x193 ;
  assign n5233 = ~x51 & n5232 ;
  assign n5234 = n5233 ^ x193 ;
  assign n5235 = ~x299 & n5234 ;
  assign n5236 = n5235 ^ x299 ;
  assign n5251 = ~x72 & n2956 ;
  assign n5252 = ~x51 & x222 ;
  assign n5253 = ~x223 & n1209 ;
  assign n5254 = n5252 & n5253 ;
  assign n5255 = ~x287 & n2655 ;
  assign n5256 = x180 & n5255 ;
  assign n5257 = n5256 ^ x224 ;
  assign n5258 = x224 & n5257 ;
  assign n5259 = n5254 & n5258 ;
  assign n5260 = n5259 ^ n5254 ;
  assign n5261 = n5251 & n5260 ;
  assign n5262 = ~n5236 & ~n5261 ;
  assign n5263 = ~n5250 & ~n5262 ;
  assign n5221 = ~x39 & ~n4386 ;
  assign n5222 = ~n5136 & n5221 ;
  assign n5223 = n1762 & n5222 ;
  assign n5224 = n5223 ^ n5221 ;
  assign n5225 = n2957 & ~n5224 ;
  assign n5237 = n5228 & n5236 ;
  assign n5188 = n5154 ^ x133 ;
  assign n5189 = n5188 ^ x125 ;
  assign n5190 = n2965 & n5189 ;
  assign n5238 = n5237 ^ n5190 ;
  assign n5239 = n5225 & ~n5238 ;
  assign n5268 = n5239 & ~n5263 ;
  assign n5269 = x39 & n5268 ;
  assign n5270 = n5269 ^ x39 ;
  assign n5240 = n5239 ^ n5238 ;
  assign n5241 = n5240 ^ x39 ;
  assign n5271 = n5270 ^ n5241 ;
  assign n5272 = ~x87 & n5271 ;
  assign n5273 = n1290 & n5272 ;
  assign n5277 = x39 & n2832 ;
  assign n5278 = n2957 & n5251 ;
  assign n5279 = n5277 & n5278 ;
  assign n5284 = n5273 & n5279 ;
  assign n5285 = ~n5263 & n5284 ;
  assign n5286 = n5285 ^ n5263 ;
  assign n5274 = n5273 ^ n1290 ;
  assign n5275 = n5274 ^ n5263 ;
  assign n5287 = n5286 ^ n5275 ;
  assign n5290 = x162 ^ x140 ;
  assign n5291 = x299 & n5290 ;
  assign n5292 = n5291 ^ x140 ;
  assign n5293 = n4926 & n5292 ;
  assign n5294 = n5287 & n5293 ;
  assign n5191 = ~n1290 & n3219 ;
  assign n5200 = n5199 ^ x162 ;
  assign n5203 = ~x87 & n5200 ;
  assign n5204 = n5203 ^ x162 ;
  assign n5205 = n5191 & n5204 ;
  assign n5206 = n5205 ^ n1290 ;
  assign n5207 = ~n5190 & ~n5206 ;
  assign n5208 = n1282 & n5139 ;
  assign n5209 = n3219 & n5208 ;
  assign n5210 = x197 ^ x145 ;
  assign n5211 = x299 & n5210 ;
  assign n5212 = n5211 ^ x145 ;
  assign n5213 = n5212 ^ n3740 ;
  assign n5216 = n5135 & n5213 ;
  assign n5217 = n5216 ^ n3740 ;
  assign n5218 = n5209 & n5217 ;
  assign n5219 = n5218 ^ n5208 ;
  assign n5220 = ~n5207 & ~n5219 ;
  assign n5289 = n5287 ^ n5220 ;
  assign n5295 = n5294 ^ n5289 ;
  assign n5296 = n2965 & ~n5208 ;
  assign n5297 = n5149 ^ x126 ;
  assign n5302 = ~x130 & n5148 ;
  assign n5303 = n5302 ^ n5150 ;
  assign n5304 = ~n5151 & n5303 ;
  assign n5305 = n5297 & ~n5304 ;
  assign n5306 = n5296 & n5305 ;
  assign n5307 = n5306 ^ n5208 ;
  assign n5308 = ~n5144 & n5307 ;
  assign n5309 = n5243 ^ n2676 ;
  assign n5315 = x182 & n5243 ;
  assign n5316 = n5315 ^ n2832 ;
  assign n5317 = n1935 & ~n5316 ;
  assign n5318 = n5317 ^ n5243 ;
  assign n5319 = ~n5309 & n5318 ;
  assign n5320 = n5317 ^ n2832 ;
  assign n5321 = n5320 ^ x160 ;
  assign n5322 = n5321 ^ n5317 ;
  assign n5323 = n5319 & ~n5322 ;
  assign n5324 = n5323 ^ n5320 ;
  assign n5325 = n2962 & n5324 ;
  assign n5326 = ~n1290 & n4927 ;
  assign n5327 = x166 ^ x153 ;
  assign n5330 = x51 & ~n5327 ;
  assign n5331 = n5330 ^ x166 ;
  assign n5332 = n5326 & ~n5331 ;
  assign n5333 = ~n2965 & ~n5332 ;
  assign n5334 = ~n5325 & ~n5333 ;
  assign n5335 = ~n5308 & n5334 ;
  assign n5354 = n4931 ^ n3810 ;
  assign n5357 = ~n5135 & n5354 ;
  assign n5358 = n5357 ^ n3810 ;
  assign n5359 = n5208 & n5358 ;
  assign n5346 = x299 ^ x185 ;
  assign n5347 = n5346 ^ x150 ;
  assign n5348 = n1537 & n5347 ;
  assign n5349 = n5348 ^ x150 ;
  assign n5341 = ~n1209 & ~n4482 ;
  assign n5336 = x175 ^ x153 ;
  assign n5337 = ~x299 & n5336 ;
  assign n5338 = n5337 ^ x153 ;
  assign n5342 = n5341 ^ n5338 ;
  assign n5343 = ~x51 & n5342 ;
  assign n5344 = n5343 ^ n5338 ;
  assign n5345 = n1290 & n5344 ;
  assign n5350 = n5349 ^ n5345 ;
  assign n5351 = ~x87 & n5350 ;
  assign n5352 = n5351 ^ n5349 ;
  assign n5360 = n5359 ^ n5352 ;
  assign n5361 = n3219 & n5360 ;
  assign n5362 = ~n5335 & ~n5361 ;
  assign n5363 = n2608 ^ x127 ;
  assign n5368 = x250 & n3250 ;
  assign n5369 = n5363 & n5368 ;
  assign n5370 = n5369 ^ n5363 ;
  assign n5371 = n5370 ^ n2608 ;
  assign n5372 = x94 & ~n5371 ;
  assign n5373 = x129 & ~n5372 ;
  assign n5374 = ~n4621 & n5373 ;
  assign n5375 = ~x250 & n3483 ;
  assign n5383 = ~n3250 & n5375 ;
  assign n5384 = ~x100 & n5383 ;
  assign n5385 = n5384 ^ x100 ;
  assign n5376 = n5375 ^ x129 ;
  assign n5377 = n5376 ^ x100 ;
  assign n5386 = n5385 ^ n5377 ;
  assign n5387 = n1275 & ~n5386 ;
  assign n5388 = ~n1341 & ~n5387 ;
  assign n5389 = ~n1919 & ~n5388 ;
  assign n5390 = ~n1290 & ~n4926 ;
  assign n5409 = n5152 ^ x130 ;
  assign n5410 = n1209 & n5409 ;
  assign n5411 = n5148 & n5410 ;
  assign n5412 = n5152 & n5411 ;
  assign n5413 = n5412 ^ n5410 ;
  assign n5414 = n5413 ^ n1209 ;
  assign n5391 = n1273 & ~n3233 ;
  assign n5395 = n2825 & n5243 ;
  assign n5400 = n5391 & n5395 ;
  assign n5401 = n5292 & n5400 ;
  assign n5402 = n5401 ^ n5292 ;
  assign n5392 = n5391 ^ n1273 ;
  assign n5393 = n5392 ^ n5292 ;
  assign n5403 = n5402 ^ n5393 ;
  assign n5404 = x39 & ~n5403 ;
  assign n5405 = n5225 & ~n5404 ;
  assign n5406 = ~x87 & n1290 ;
  assign n5407 = ~n5405 & n5406 ;
  assign n5408 = ~n5279 & n5407 ;
  assign n5415 = n5408 & n5414 ;
  assign n5416 = n5415 ^ n5407 ;
  assign n5417 = ~n1209 & n5416 ;
  assign n5418 = n3529 & n5417 ;
  assign n5419 = n5418 ^ n5416 ;
  assign n5420 = ~n5414 & ~n5419 ;
  assign n5421 = n5390 & n5420 ;
  assign n5425 = ~n1209 & n3219 ;
  assign n5430 = n5421 & n5425 ;
  assign n5431 = x169 & n5430 ;
  assign n5432 = n5431 ^ x169 ;
  assign n5422 = n5421 ^ n5419 ;
  assign n5423 = n5422 ^ x169 ;
  assign n5433 = n5432 ^ n5423 ;
  assign n5434 = ~x51 & n5433 ;
  assign n5437 = n1537 & n3760 ;
  assign n5438 = n5437 ^ x167 ;
  assign n5439 = n4926 & n5438 ;
  assign n5440 = n5439 ^ x87 ;
  assign n5441 = ~n5434 & ~n5440 ;
  assign n5442 = n2832 & n2962 ;
  assign n5443 = n2965 & ~n5442 ;
  assign n5444 = ~n5139 & n5443 ;
  assign n5445 = n3219 & n4470 ;
  assign n5446 = n5133 & n5445 ;
  assign n5447 = n5446 ^ n5133 ;
  assign n5449 = x183 & n1420 ;
  assign n5448 = x149 & n2674 ;
  assign n5450 = n5449 ^ n5448 ;
  assign n5451 = ~n5447 & n5450 ;
  assign n5452 = n5243 & n5451 ;
  assign n5453 = n2965 & n5452 ;
  assign n5454 = ~n5444 & ~n5453 ;
  assign n5455 = x132 ^ x126 ;
  assign n5456 = n5455 ^ n5304 ;
  assign n5457 = n5456 ^ x132 ;
  assign n5460 = n5149 & ~n5457 ;
  assign n5461 = n5460 ^ x132 ;
  assign n5462 = ~n5144 & n5461 ;
  assign n5463 = ~n5454 & ~n5462 ;
  assign n5464 = x190 ^ x168 ;
  assign n5467 = ~n1537 & n5464 ;
  assign n5468 = n5467 ^ x190 ;
  assign n5469 = n5114 & n5468 ;
  assign n5470 = n5469 ^ n2964 ;
  assign n5474 = ~n1290 & n3532 ;
  assign n5475 = n5474 ^ n3533 ;
  assign n5476 = n4926 & ~n5475 ;
  assign n5477 = n5476 ^ n3219 ;
  assign n5478 = n2963 & n5477 ;
  assign n5481 = n1537 & n4978 ;
  assign n5482 = n5481 ^ x151 ;
  assign n5483 = n5478 & ~n5482 ;
  assign n5484 = n5483 ^ n5477 ;
  assign n5485 = n5470 & n5484 ;
  assign n5486 = ~n5463 & ~n5485 ;
  assign n5487 = n5208 & ~n5447 ;
  assign n5488 = n5486 & n5487 ;
  assign n5489 = n5488 ^ n5486 ;
  assign n5490 = x183 ^ x149 ;
  assign n5493 = ~n1537 & n5490 ;
  assign n5494 = n5493 ^ x183 ;
  assign n5495 = n4926 & n5494 ;
  assign n5506 = n5188 & ~n5495 ;
  assign n5507 = n5443 & n5506 ;
  assign n5508 = n5507 ^ n5443 ;
  assign n5496 = ~x86 & n3456 ;
  assign n5497 = ~n3562 & n5496 ;
  assign n5498 = n5497 ^ n3562 ;
  assign n5499 = n5498 ^ n5495 ;
  assign n5500 = n5499 ^ n5443 ;
  assign n5509 = n5508 ^ n5500 ;
  assign n5510 = ~n5208 & n5509 ;
  assign n5511 = n5510 ^ n5498 ;
  assign n5512 = ~x72 & ~n3233 ;
  assign n5513 = n5140 & n5512 ;
  assign n5521 = n5395 & n5513 ;
  assign n5522 = n5212 & n5521 ;
  assign n5523 = n5522 ^ n5212 ;
  assign n5514 = n5513 ^ n5140 ;
  assign n5515 = n5514 ^ n5212 ;
  assign n5524 = n5523 ^ n5515 ;
  assign n5525 = ~n4621 & n5524 ;
  assign n5526 = ~n5511 & ~n5525 ;
  assign n5527 = ~n2964 & ~n5139 ;
  assign n5551 = x192 ^ x171 ;
  assign n5554 = ~n1537 & n5551 ;
  assign n5555 = n5554 ^ x192 ;
  assign n5556 = n3219 & n5555 ;
  assign n5528 = ~x136 & n5153 ;
  assign n5534 = ~x135 & n5528 ;
  assign n5529 = n5154 ^ x134 ;
  assign n5535 = n5534 ^ n5529 ;
  assign n5536 = ~n5144 & ~n5535 ;
  assign n5537 = n5536 ^ n5512 ;
  assign n5538 = n5141 & n5537 ;
  assign n5546 = n3533 & n5538 ;
  assign n5547 = n5395 & n5546 ;
  assign n5548 = n5547 ^ n5395 ;
  assign n5539 = n5538 ^ n5141 ;
  assign n5540 = n5539 ^ n5395 ;
  assign n5549 = n5548 ^ n5540 ;
  assign n5550 = ~n5536 & ~n5549 ;
  assign n5557 = n5556 ^ n5550 ;
  assign n5558 = ~n1209 & ~n5557 ;
  assign n5559 = n5558 ^ n5550 ;
  assign n5560 = n5527 & n5559 ;
  assign n5573 = x194 ^ x170 ;
  assign n5576 = n1537 & n5573 ;
  assign n5577 = n5576 ^ x170 ;
  assign n5578 = n5425 & n5577 ;
  assign n5562 = x185 & n1420 ;
  assign n5561 = x150 & n2674 ;
  assign n5563 = n5562 ^ n5561 ;
  assign n5564 = n5243 & n5563 ;
  assign n5565 = n5442 & ~n5564 ;
  assign n5566 = n1209 & ~n5565 ;
  assign n5567 = ~n5144 & n5566 ;
  assign n5568 = n5528 ^ n5154 ;
  assign n5569 = n5568 ^ x135 ;
  assign n5570 = n5567 & n5569 ;
  assign n5571 = n5570 ^ n5566 ;
  assign n5579 = n5578 ^ n5571 ;
  assign n5580 = n5527 & ~n5579 ;
  assign n5587 = n5153 ^ x136 ;
  assign n5588 = n1209 & ~n5148 ;
  assign n5589 = n5587 & n5588 ;
  assign n5583 = n1537 & n3766 ;
  assign n5584 = n5583 ^ x148 ;
  assign n5585 = n5425 & n5584 ;
  assign n5586 = n5585 ^ n1209 ;
  assign n5590 = n5589 ^ n5586 ;
  assign n5591 = ~n5442 & n5590 ;
  assign n5592 = ~n2964 & ~n5591 ;
  assign n5593 = n2958 & ~n5224 ;
  assign n5601 = n3219 & n3768 ;
  assign n5595 = x184 & n1420 ;
  assign n5594 = x163 & n2674 ;
  assign n5596 = n5595 ^ n5594 ;
  assign n5597 = n5243 & n5596 ;
  assign n5598 = ~n3233 & ~n5597 ;
  assign n5599 = n5251 & ~n5598 ;
  assign n5600 = x39 & ~n5599 ;
  assign n5602 = n5601 ^ n5600 ;
  assign n5603 = n1209 & ~n5602 ;
  assign n5604 = n5603 ^ n5601 ;
  assign n5605 = n5593 & n5604 ;
  assign n5606 = n5592 & ~n5605 ;
  assign n5608 = ~x210 & n4046 ;
  assign n5607 = ~x198 & n4052 ;
  assign n5609 = n5608 ^ n5607 ;
  assign n5610 = n4070 & n5609 ;
  assign n5611 = n3219 & n5610 ;
  assign n5612 = n5611 ^ x137 ;
  assign n5613 = x39 & n5612 ;
  assign n5614 = n5613 ^ x137 ;
  assign n5615 = n1289 & n3210 ;
  assign n5620 = n2689 & n3537 ;
  assign n5621 = n5620 ^ n3625 ;
  assign n5622 = x39 & n5621 ;
  assign n5623 = n5622 ^ n3625 ;
  assign n5624 = n5615 & n5623 ;
  assign n5625 = n3703 & ~n5624 ;
  assign n5626 = n1340 & n5625 ;
  assign n5632 = ~x195 & ~x196 ;
  assign n5633 = n5632 ^ n3545 ;
  assign n5634 = ~n3546 & n5633 ;
  assign n5627 = x139 ^ x138 ;
  assign n5635 = n5634 ^ n5627 ;
  assign n5636 = n5635 ^ x138 ;
  assign n5639 = n3544 & ~n5636 ;
  assign n5640 = n5639 ^ x138 ;
  assign n5641 = n5626 & n5640 ;
  assign n5642 = n5641 ^ n5601 ;
  assign n5643 = ~n4402 & ~n5642 ;
  assign n5644 = n5643 ^ n5601 ;
  assign n5645 = n3549 ^ n3544 ;
  assign n5646 = n5645 ^ x139 ;
  assign n5647 = n5626 & n5646 ;
  assign n5648 = n5647 ^ n3529 ;
  assign n5649 = n4402 & ~n5648 ;
  assign n5650 = n5649 ^ n5647 ;
  assign n5727 = n3237 ^ n2966 ;
  assign n5671 = n4346 ^ n3237 ;
  assign n5728 = n5727 ^ n5671 ;
  assign n5652 = ~x120 & ~x287 ;
  assign n5653 = n3970 & n5652 ;
  assign n5654 = n5653 ^ x120 ;
  assign n5732 = n5728 ^ n5654 ;
  assign n5730 = n5728 ^ n2708 ;
  assign n5731 = n5730 ^ n5671 ;
  assign n5735 = n5732 ^ n5731 ;
  assign n5736 = n5735 ^ n5727 ;
  assign n5737 = n5736 ^ n3237 ;
  assign n5651 = n2966 ^ n2708 ;
  assign n5655 = n5654 ^ n5651 ;
  assign n5710 = n5727 ^ n5655 ;
  assign n5711 = n5710 ^ n5671 ;
  assign n5712 = n5730 ^ n5711 ;
  assign n5689 = n4346 & ~n5671 ;
  assign n5690 = n5710 ^ n5689 ;
  assign n5670 = n3237 ^ n2708 ;
  assign n5691 = n5690 ^ n5670 ;
  assign n5692 = n5691 ^ n3237 ;
  assign n5695 = ~n5655 & n5692 ;
  assign n5698 = n5736 ^ n5710 ;
  assign n5699 = n5737 ^ n5698 ;
  assign n5700 = n5651 & n5699 ;
  assign n5701 = n5695 & n5700 ;
  assign n5702 = n5701 ^ n5689 ;
  assign n5703 = n5712 ^ n5702 ;
  assign n5672 = n5671 ^ n5670 ;
  assign n5726 = n5703 ^ n5672 ;
  assign n5738 = n5737 ^ n5726 ;
  assign n5739 = ~x841 & n1266 ;
  assign n5744 = n1557 & n5739 ;
  assign n5740 = ~x45 & ~x47 ;
  assign n5741 = ~x102 & ~n3952 ;
  assign n5742 = n5740 & n5741 ;
  assign n5745 = n5744 ^ n5742 ;
  assign n5746 = ~x252 & ~n5745 ;
  assign n5754 = ~x47 & n5746 ;
  assign n5755 = ~n1244 & n5754 ;
  assign n5756 = n5755 ^ n1244 ;
  assign n5747 = n5746 ^ n5745 ;
  assign n5748 = n5747 ^ n1244 ;
  assign n5757 = n5756 ^ n5748 ;
  assign n5758 = ~x40 & n5757 ;
  assign n5759 = ~n4381 & n5758 ;
  assign n5760 = ~n4621 & n5759 ;
  assign n5762 = ~n2698 & n3984 ;
  assign n5763 = n5760 & n5762 ;
  assign n5761 = n5760 ^ n4621 ;
  assign n5764 = n5763 ^ n5761 ;
  assign n5765 = ~n5738 & n5764 ;
  assign n5766 = n3009 & ~n5765 ;
  assign n5767 = x832 & n3009 ;
  assign n5768 = ~n5766 & ~n5767 ;
  assign n5844 = x761 ^ x140 ;
  assign n5769 = x621 & x1091 ;
  assign n5770 = x1156 ^ x629 ;
  assign n5771 = x1153 ^ x608 ;
  assign n5772 = x1159 ^ x619 ;
  assign n5773 = x1160 ^ x644 ;
  assign n5774 = x1158 ^ x626 ;
  assign n5782 = x1157 ^ x630 ;
  assign n5775 = x1155 ^ x609 ;
  assign n5776 = x1154 ^ x618 ;
  assign n5777 = x781 & n5776 ;
  assign n5778 = x603 & ~n5777 ;
  assign n5779 = x785 & n5778 ;
  assign n5780 = n5775 & n5779 ;
  assign n5781 = n5780 ^ n5778 ;
  assign n5783 = x787 & n5781 ;
  assign n5784 = n5782 & n5783 ;
  assign n5785 = n5784 ^ n5781 ;
  assign n5786 = x788 & n5785 ;
  assign n5787 = n5774 & n5786 ;
  assign n5788 = n5787 ^ n5785 ;
  assign n5789 = x790 & n5788 ;
  assign n5790 = n5773 & n5789 ;
  assign n5791 = n5790 ^ n5788 ;
  assign n5792 = x789 & n5791 ;
  assign n5793 = n5772 & n5792 ;
  assign n5794 = n5793 ^ n5791 ;
  assign n5795 = x778 & n5794 ;
  assign n5796 = n5771 & n5795 ;
  assign n5797 = n5796 ^ n5794 ;
  assign n5798 = x792 & n5797 ;
  assign n5799 = n5770 & n5798 ;
  assign n5800 = n5799 ^ n5797 ;
  assign n5801 = n5769 & n5800 ;
  assign n5802 = n5801 ^ n5800 ;
  assign n5805 = x665 & x1091 ;
  assign n5806 = x1159 ^ x648 ;
  assign n5807 = x1156 ^ x628 ;
  assign n5808 = x1157 ^ x647 ;
  assign n5809 = x1154 ^ x627 ;
  assign n5821 = x1155 ^ x660 ;
  assign n5810 = x1153 ^ x625 ;
  assign n5811 = x1158 ^ x641 ;
  assign n5812 = x1160 ^ x715 ;
  assign n5813 = x790 & n5812 ;
  assign n5814 = x788 & ~n5813 ;
  assign n5815 = n5811 & n5814 ;
  assign n5816 = n5815 ^ n5813 ;
  assign n5817 = x680 & ~n5816 ;
  assign n5818 = x778 & n5817 ;
  assign n5819 = n5810 & n5818 ;
  assign n5820 = n5819 ^ n5817 ;
  assign n5822 = x785 & n5820 ;
  assign n5823 = n5821 & n5822 ;
  assign n5824 = n5823 ^ n5820 ;
  assign n5825 = x781 & n5824 ;
  assign n5826 = n5809 & n5825 ;
  assign n5827 = n5826 ^ n5824 ;
  assign n5828 = x787 & n5827 ;
  assign n5829 = n5808 & n5828 ;
  assign n5830 = n5829 ^ n5827 ;
  assign n5831 = x792 & n5830 ;
  assign n5832 = n5807 & n5831 ;
  assign n5833 = n5832 ^ n5830 ;
  assign n5834 = x789 & n5833 ;
  assign n5835 = n5806 & n5834 ;
  assign n5836 = n5835 ^ n5833 ;
  assign n5837 = n5805 & n5836 ;
  assign n5838 = n5837 ^ n5836 ;
  assign n5841 = ~x738 & n5838 ;
  assign n5842 = n5841 ^ x761 ;
  assign n5843 = ~n5802 & ~n5842 ;
  assign n5845 = n5844 ^ n5843 ;
  assign n5846 = ~n5768 & n5845 ;
  assign n5847 = n5846 ^ x140 ;
  assign n5855 = x749 ^ x141 ;
  assign n5852 = x706 & n5838 ;
  assign n5853 = n5852 ^ x749 ;
  assign n5854 = ~n5802 & n5853 ;
  assign n5856 = n5855 ^ n5854 ;
  assign n5857 = ~n5768 & ~n5856 ;
  assign n5858 = n5857 ^ x141 ;
  assign n5866 = x743 ^ x142 ;
  assign n5863 = x735 & n5838 ;
  assign n5864 = n5863 ^ x743 ;
  assign n5865 = ~n5802 & n5864 ;
  assign n5867 = n5866 ^ n5865 ;
  assign n5868 = ~n5768 & n5867 ;
  assign n5869 = n5868 ^ x142 ;
  assign n5877 = x774 ^ x143 ;
  assign n5874 = x687 & n5838 ;
  assign n5875 = n5874 ^ x774 ;
  assign n5876 = ~n5802 & ~n5875 ;
  assign n5878 = n5877 ^ n5876 ;
  assign n5879 = ~n5768 & n5878 ;
  assign n5880 = n5879 ^ x143 ;
  assign n5888 = x758 ^ x144 ;
  assign n5885 = x736 & n5838 ;
  assign n5886 = n5885 ^ x758 ;
  assign n5887 = ~n5802 & n5886 ;
  assign n5889 = n5888 ^ n5887 ;
  assign n5890 = ~n5768 & n5889 ;
  assign n5891 = n5890 ^ x144 ;
  assign n5899 = x767 ^ x145 ;
  assign n5896 = ~x698 & n5838 ;
  assign n5897 = n5896 ^ x767 ;
  assign n5898 = ~n5802 & ~n5897 ;
  assign n5900 = n5899 ^ n5898 ;
  assign n5901 = ~n5768 & n5900 ;
  assign n5902 = n5901 ^ x145 ;
  assign n5908 = x743 ^ x146 ;
  assign n5905 = x735 & x907 ;
  assign n5906 = n5905 ^ x743 ;
  assign n5907 = ~x947 & n5906 ;
  assign n5909 = n5908 ^ n5907 ;
  assign n5910 = ~n5768 & n5909 ;
  assign n5911 = n5910 ^ x146 ;
  assign n5919 = x770 ^ x147 ;
  assign n5916 = x726 & x907 ;
  assign n5917 = n5916 ^ x770 ;
  assign n5918 = ~x947 & ~n5917 ;
  assign n5920 = n5919 ^ n5918 ;
  assign n5921 = ~n5768 & n5920 ;
  assign n5922 = n5921 ^ x147 ;
  assign n5928 = x749 ^ x148 ;
  assign n5925 = x706 & x907 ;
  assign n5926 = n5925 ^ x749 ;
  assign n5927 = ~x947 & n5926 ;
  assign n5929 = n5928 ^ n5927 ;
  assign n5930 = ~n5768 & ~n5929 ;
  assign n5931 = n5930 ^ x148 ;
  assign n5954 = ~x149 & n5768 ;
  assign n5933 = n1510 & n2704 ;
  assign n5935 = n5933 ^ n2706 ;
  assign n5932 = n3234 & n3600 ;
  assign n5936 = n5933 ^ n5932 ;
  assign n5937 = n2966 & ~n5936 ;
  assign n5938 = n5654 & n5937 ;
  assign n5939 = ~n5935 & n5938 ;
  assign n5940 = n5939 ^ n5937 ;
  assign n5941 = n5940 ^ n2966 ;
  assign n5942 = n5764 & ~n5941 ;
  assign n5943 = n3009 & ~n5942 ;
  assign n5944 = ~n5767 & ~n5943 ;
  assign n5949 = ~x725 & x907 ;
  assign n5950 = n5949 ^ x755 ;
  assign n5951 = ~x947 & ~n5950 ;
  assign n5952 = n5951 ^ x755 ;
  assign n5953 = ~n5944 & ~n5952 ;
  assign n5956 = n5954 ^ n5953 ;
  assign n5966 = ~x150 & n5768 ;
  assign n5961 = ~x701 & x907 ;
  assign n5962 = n5961 ^ x751 ;
  assign n5963 = ~x947 & ~n5962 ;
  assign n5964 = n5963 ^ x751 ;
  assign n5965 = ~n5944 & ~n5964 ;
  assign n5968 = n5966 ^ n5965 ;
  assign n5976 = x745 ^ x151 ;
  assign n5973 = ~x723 & x907 ;
  assign n5974 = n5973 ^ x745 ;
  assign n5975 = ~x947 & ~n5974 ;
  assign n5977 = n5976 ^ n5975 ;
  assign n5978 = ~n5768 & n5977 ;
  assign n5979 = n5978 ^ x151 ;
  assign n5987 = x759 ^ x152 ;
  assign n5984 = x696 & x907 ;
  assign n5985 = n5984 ^ x759 ;
  assign n5986 = ~x947 & n5985 ;
  assign n5988 = n5987 ^ n5986 ;
  assign n5989 = ~n5768 & n5988 ;
  assign n5990 = n5989 ^ x152 ;
  assign n5998 = x766 ^ x153 ;
  assign n5995 = x700 & x907 ;
  assign n5996 = n5995 ^ x766 ;
  assign n5997 = ~x947 & n5996 ;
  assign n5999 = n5998 ^ n5997 ;
  assign n6000 = ~n5768 & ~n5999 ;
  assign n6001 = n6000 ^ x153 ;
  assign n6011 = ~x154 & n5768 ;
  assign n6006 = ~x704 & x907 ;
  assign n6007 = n6006 ^ x742 ;
  assign n6008 = ~x947 & ~n6007 ;
  assign n6009 = n6008 ^ x742 ;
  assign n6010 = ~n5944 & ~n6009 ;
  assign n6013 = n6011 ^ n6010 ;
  assign n6023 = ~x155 & n5768 ;
  assign n6018 = ~x686 & x907 ;
  assign n6019 = n6018 ^ x757 ;
  assign n6020 = ~x947 & ~n6019 ;
  assign n6021 = n6020 ^ x757 ;
  assign n6022 = ~n5944 & ~n6021 ;
  assign n6025 = n6023 ^ n6022 ;
  assign n6035 = ~x156 & n5768 ;
  assign n6030 = ~x724 & x907 ;
  assign n6031 = n6030 ^ x741 ;
  assign n6032 = ~x947 & ~n6031 ;
  assign n6033 = n6032 ^ x741 ;
  assign n6034 = ~n5944 & ~n6033 ;
  assign n6037 = n6035 ^ n6034 ;
  assign n6045 = x760 ^ x157 ;
  assign n6042 = ~x688 & x907 ;
  assign n6043 = n6042 ^ x760 ;
  assign n6044 = ~x947 & ~n6043 ;
  assign n6046 = n6045 ^ n6044 ;
  assign n6047 = ~n5768 & n6046 ;
  assign n6048 = n6047 ^ x157 ;
  assign n6058 = ~x158 & n5768 ;
  assign n6053 = ~x702 & x907 ;
  assign n6054 = n6053 ^ x753 ;
  assign n6055 = ~x947 & ~n6054 ;
  assign n6056 = n6055 ^ x753 ;
  assign n6057 = ~n5944 & ~n6056 ;
  assign n6060 = n6058 ^ n6057 ;
  assign n6068 = x754 ^ x159 ;
  assign n6065 = ~x709 & x907 ;
  assign n6066 = n6065 ^ x754 ;
  assign n6067 = ~x947 & ~n6066 ;
  assign n6069 = n6068 ^ n6067 ;
  assign n6070 = ~n5768 & n6069 ;
  assign n6071 = n6070 ^ x159 ;
  assign n6079 = x756 ^ x160 ;
  assign n6076 = ~x734 & x907 ;
  assign n6077 = n6076 ^ x756 ;
  assign n6078 = ~x947 & ~n6077 ;
  assign n6080 = n6079 ^ n6078 ;
  assign n6081 = ~n5768 & n6080 ;
  assign n6082 = n6081 ^ x160 ;
  assign n6088 = x758 ^ x161 ;
  assign n6085 = x736 & x907 ;
  assign n6086 = n6085 ^ x758 ;
  assign n6087 = ~x947 & n6086 ;
  assign n6089 = n6088 ^ n6087 ;
  assign n6090 = ~n5768 & n6089 ;
  assign n6091 = n6090 ^ x161 ;
  assign n6097 = x761 ^ x162 ;
  assign n6094 = ~x738 & x907 ;
  assign n6095 = n6094 ^ x761 ;
  assign n6096 = ~x947 & ~n6095 ;
  assign n6098 = n6097 ^ n6096 ;
  assign n6099 = ~n5768 & n6098 ;
  assign n6100 = n6099 ^ x162 ;
  assign n6108 = x777 ^ x163 ;
  assign n6105 = ~x737 & x907 ;
  assign n6106 = n6105 ^ x777 ;
  assign n6107 = ~x947 & ~n6106 ;
  assign n6109 = n6108 ^ n6107 ;
  assign n6110 = ~n5768 & n6109 ;
  assign n6111 = n6110 ^ x163 ;
  assign n6119 = x752 ^ x164 ;
  assign n6116 = x703 & x907 ;
  assign n6117 = n6116 ^ x752 ;
  assign n6118 = ~x947 & ~n6117 ;
  assign n6120 = n6119 ^ n6118 ;
  assign n6121 = ~n5768 & n6120 ;
  assign n6122 = n6121 ^ x164 ;
  assign n6130 = ~x165 & n5768 ;
  assign n6125 = x687 & x907 ;
  assign n6126 = n6125 ^ x774 ;
  assign n6127 = ~x947 & ~n6126 ;
  assign n6128 = n6127 ^ x774 ;
  assign n6129 = ~n5944 & ~n6128 ;
  assign n6132 = n6130 ^ n6129 ;
  assign n6140 = x772 ^ x166 ;
  assign n6137 = x727 & x907 ;
  assign n6138 = n6137 ^ x772 ;
  assign n6139 = ~x947 & n6138 ;
  assign n6141 = n6140 ^ n6139 ;
  assign n6142 = ~n5768 & n6141 ;
  assign n6143 = n6142 ^ x166 ;
  assign n6151 = x768 ^ x167 ;
  assign n6148 = x705 & x907 ;
  assign n6149 = n6148 ^ x768 ;
  assign n6150 = ~x947 & ~n6149 ;
  assign n6152 = n6151 ^ n6150 ;
  assign n6153 = ~n5768 & n6152 ;
  assign n6154 = n6153 ^ x167 ;
  assign n6162 = x763 ^ x168 ;
  assign n6159 = x699 & x907 ;
  assign n6160 = n6159 ^ x763 ;
  assign n6161 = ~x947 & n6160 ;
  assign n6163 = n6162 ^ n6161 ;
  assign n6164 = ~n5768 & ~n6163 ;
  assign n6165 = n6164 ^ x168 ;
  assign n6173 = x746 ^ x169 ;
  assign n6170 = x729 & x907 ;
  assign n6171 = n6170 ^ x746 ;
  assign n6172 = ~x947 & n6171 ;
  assign n6174 = n6173 ^ n6172 ;
  assign n6175 = ~n5768 & ~n6174 ;
  assign n6176 = n6175 ^ x169 ;
  assign n6184 = x748 ^ x170 ;
  assign n6181 = x730 & x907 ;
  assign n6182 = n6181 ^ x748 ;
  assign n6183 = ~x947 & n6182 ;
  assign n6185 = n6184 ^ n6183 ;
  assign n6186 = ~n5768 & ~n6185 ;
  assign n6187 = n6186 ^ x170 ;
  assign n6195 = x764 ^ x171 ;
  assign n6192 = x691 & x907 ;
  assign n6193 = n6192 ^ x764 ;
  assign n6194 = ~x947 & n6193 ;
  assign n6196 = n6195 ^ n6194 ;
  assign n6197 = ~n5768 & ~n6196 ;
  assign n6198 = n6197 ^ x171 ;
  assign n6206 = x739 ^ x172 ;
  assign n6203 = x690 & x907 ;
  assign n6204 = n6203 ^ x739 ;
  assign n6205 = ~x947 & n6204 ;
  assign n6207 = n6206 ^ n6205 ;
  assign n6208 = ~n5768 & ~n6207 ;
  assign n6209 = n6208 ^ x172 ;
  assign n6215 = x745 ^ x173 ;
  assign n6212 = ~x723 & n5838 ;
  assign n6213 = n6212 ^ x745 ;
  assign n6214 = ~n5802 & ~n6213 ;
  assign n6216 = n6215 ^ n6214 ;
  assign n6217 = ~n5768 & n6216 ;
  assign n6218 = n6217 ^ x173 ;
  assign n6224 = x759 ^ x174 ;
  assign n6221 = x696 & n5838 ;
  assign n6222 = n6221 ^ x759 ;
  assign n6223 = ~n5802 & n6222 ;
  assign n6225 = n6224 ^ n6223 ;
  assign n6226 = ~n5768 & n6225 ;
  assign n6227 = n6226 ^ x174 ;
  assign n6233 = x766 ^ x175 ;
  assign n6230 = x700 & n5838 ;
  assign n6231 = n6230 ^ x766 ;
  assign n6232 = ~n5802 & n6231 ;
  assign n6234 = n6233 ^ n6232 ;
  assign n6235 = ~n5768 & ~n6234 ;
  assign n6236 = n6235 ^ x175 ;
  assign n6242 = x742 ^ x176 ;
  assign n6239 = ~x704 & n5838 ;
  assign n6240 = n6239 ^ x742 ;
  assign n6241 = ~n5802 & ~n6240 ;
  assign n6243 = n6242 ^ n6241 ;
  assign n6244 = ~n5768 & n6243 ;
  assign n6245 = n6244 ^ x176 ;
  assign n6251 = x757 ^ x177 ;
  assign n6248 = ~x686 & n5838 ;
  assign n6249 = n6248 ^ x757 ;
  assign n6250 = ~n5802 & ~n6249 ;
  assign n6252 = n6251 ^ n6250 ;
  assign n6253 = ~n5768 & n6252 ;
  assign n6254 = n6253 ^ x177 ;
  assign n6260 = x760 ^ x178 ;
  assign n6257 = ~x688 & n5838 ;
  assign n6258 = n6257 ^ x760 ;
  assign n6259 = ~n5802 & ~n6258 ;
  assign n6261 = n6260 ^ n6259 ;
  assign n6262 = ~n5768 & n6261 ;
  assign n6263 = n6262 ^ x178 ;
  assign n6269 = x741 ^ x179 ;
  assign n6266 = ~x724 & n5838 ;
  assign n6267 = n6266 ^ x741 ;
  assign n6268 = ~n5802 & ~n6267 ;
  assign n6270 = n6269 ^ n6268 ;
  assign n6271 = ~n5768 & n6270 ;
  assign n6272 = n6271 ^ x179 ;
  assign n6278 = x753 ^ x180 ;
  assign n6275 = ~x702 & n5838 ;
  assign n6276 = n6275 ^ x753 ;
  assign n6277 = ~n5802 & ~n6276 ;
  assign n6279 = n6278 ^ n6277 ;
  assign n6280 = ~n5768 & n6279 ;
  assign n6281 = n6280 ^ x180 ;
  assign n6287 = x754 ^ x181 ;
  assign n6284 = ~x709 & n5838 ;
  assign n6285 = n6284 ^ x754 ;
  assign n6286 = ~n5802 & ~n6285 ;
  assign n6288 = n6287 ^ n6286 ;
  assign n6289 = ~n5768 & n6288 ;
  assign n6290 = n6289 ^ x181 ;
  assign n6296 = x756 ^ x182 ;
  assign n6293 = ~x734 & n5838 ;
  assign n6294 = n6293 ^ x756 ;
  assign n6295 = ~n5802 & ~n6294 ;
  assign n6297 = n6296 ^ n6295 ;
  assign n6298 = ~n5768 & n6297 ;
  assign n6299 = n6298 ^ x182 ;
  assign n6305 = x755 ^ x183 ;
  assign n6302 = ~x725 & n5838 ;
  assign n6303 = n6302 ^ x755 ;
  assign n6304 = ~n5802 & ~n6303 ;
  assign n6306 = n6305 ^ n6304 ;
  assign n6307 = ~n5768 & n6306 ;
  assign n6308 = n6307 ^ x183 ;
  assign n6314 = x777 ^ x184 ;
  assign n6311 = ~x737 & n5838 ;
  assign n6312 = n6311 ^ x777 ;
  assign n6313 = ~n5802 & ~n6312 ;
  assign n6315 = n6314 ^ n6313 ;
  assign n6316 = ~n5768 & n6315 ;
  assign n6317 = n6316 ^ x184 ;
  assign n6323 = x751 ^ x185 ;
  assign n6320 = ~x701 & n5838 ;
  assign n6321 = n6320 ^ x751 ;
  assign n6322 = ~n5802 & ~n6321 ;
  assign n6324 = n6323 ^ n6322 ;
  assign n6325 = ~n5768 & n6324 ;
  assign n6326 = n6325 ^ x185 ;
  assign n6332 = x752 ^ x186 ;
  assign n6329 = x703 & n5838 ;
  assign n6330 = n6329 ^ x752 ;
  assign n6331 = ~n5802 & ~n6330 ;
  assign n6333 = n6332 ^ n6331 ;
  assign n6334 = ~n5768 & n6333 ;
  assign n6335 = n6334 ^ x186 ;
  assign n6341 = x770 ^ x187 ;
  assign n6338 = x726 & n5838 ;
  assign n6339 = n6338 ^ x770 ;
  assign n6340 = ~n5802 & ~n6339 ;
  assign n6342 = n6341 ^ n6340 ;
  assign n6343 = ~n5768 & n6342 ;
  assign n6344 = n6343 ^ x187 ;
  assign n6350 = x768 ^ x188 ;
  assign n6347 = x705 & n5838 ;
  assign n6348 = n6347 ^ x768 ;
  assign n6349 = ~n5802 & ~n6348 ;
  assign n6351 = n6350 ^ n6349 ;
  assign n6352 = ~n5768 & n6351 ;
  assign n6353 = n6352 ^ x188 ;
  assign n6359 = x772 ^ x189 ;
  assign n6356 = x727 & n5838 ;
  assign n6357 = n6356 ^ x772 ;
  assign n6358 = ~n5802 & n6357 ;
  assign n6360 = n6359 ^ n6358 ;
  assign n6361 = ~n5768 & n6360 ;
  assign n6362 = n6361 ^ x189 ;
  assign n6368 = x763 ^ x190 ;
  assign n6365 = x699 & n5838 ;
  assign n6366 = n6365 ^ x763 ;
  assign n6367 = ~n5802 & n6366 ;
  assign n6369 = n6368 ^ n6367 ;
  assign n6370 = ~n5768 & ~n6369 ;
  assign n6371 = n6370 ^ x190 ;
  assign n6377 = x746 ^ x191 ;
  assign n6374 = x729 & n5838 ;
  assign n6375 = n6374 ^ x746 ;
  assign n6376 = ~n5802 & n6375 ;
  assign n6378 = n6377 ^ n6376 ;
  assign n6379 = ~n5768 & ~n6378 ;
  assign n6380 = n6379 ^ x191 ;
  assign n6386 = x764 ^ x192 ;
  assign n6383 = x691 & n5838 ;
  assign n6384 = n6383 ^ x764 ;
  assign n6385 = ~n5802 & n6384 ;
  assign n6387 = n6386 ^ n6385 ;
  assign n6388 = ~n5768 & ~n6387 ;
  assign n6389 = n6388 ^ x192 ;
  assign n6395 = x739 ^ x193 ;
  assign n6392 = x690 & n5838 ;
  assign n6393 = n6392 ^ x739 ;
  assign n6394 = ~n5802 & n6393 ;
  assign n6396 = n6395 ^ n6394 ;
  assign n6397 = ~n5768 & ~n6396 ;
  assign n6398 = n6397 ^ x193 ;
  assign n6404 = x748 ^ x194 ;
  assign n6401 = x730 & n5838 ;
  assign n6402 = n6401 ^ x748 ;
  assign n6403 = ~n5802 & n6402 ;
  assign n6405 = n6404 ^ n6403 ;
  assign n6406 = ~n5768 & ~n6405 ;
  assign n6407 = n6406 ^ x194 ;
  assign n6415 = n3548 ^ x195 ;
  assign n6416 = n6415 ^ n3549 ;
  assign n6421 = ~n5626 & n6416 ;
  assign n6412 = ~x299 & n5551 ;
  assign n6413 = n6412 ^ x171 ;
  assign n6414 = n3219 & n6413 ;
  assign n6417 = n6416 ^ n6414 ;
  assign n6422 = n6421 ^ n6417 ;
  assign n6423 = ~n4402 & ~n6422 ;
  assign n6424 = n6423 ^ n6414 ;
  assign n6430 = n3549 ^ n3547 ;
  assign n6431 = n6430 ^ x196 ;
  assign n6432 = n5626 & n6431 ;
  assign n6427 = x299 & n5573 ;
  assign n6428 = n6427 ^ x194 ;
  assign n6429 = n3219 & n6428 ;
  assign n6433 = n6432 ^ n6429 ;
  assign n6434 = n4402 & ~n6433 ;
  assign n6435 = n6434 ^ n6432 ;
  assign n6441 = x767 ^ x197 ;
  assign n6438 = ~x698 & x907 ;
  assign n6439 = n6438 ^ x767 ;
  assign n6440 = ~x947 & ~n6439 ;
  assign n6442 = n6441 ^ n6440 ;
  assign n6443 = ~n5768 & n6442 ;
  assign n6444 = n6443 ^ x197 ;
  assign n6452 = x633 ^ x198 ;
  assign n6449 = x634 & n5838 ;
  assign n6450 = n6449 ^ x633 ;
  assign n6451 = ~n5802 & n6450 ;
  assign n6453 = n6452 ^ n6451 ;
  assign n6454 = n5766 & n6453 ;
  assign n6455 = n6454 ^ x198 ;
  assign n6463 = x617 ^ x199 ;
  assign n6460 = x637 & n5838 ;
  assign n6461 = n6460 ^ x617 ;
  assign n6462 = ~n5802 & n6461 ;
  assign n6464 = n6463 ^ n6462 ;
  assign n6465 = n5766 & n6464 ;
  assign n6466 = n6465 ^ x199 ;
  assign n6474 = x606 ^ x200 ;
  assign n6471 = x643 & n5838 ;
  assign n6472 = n6471 ^ x606 ;
  assign n6473 = ~n5802 & n6472 ;
  assign n6475 = n6474 ^ n6473 ;
  assign n6476 = n5766 & n6475 ;
  assign n6477 = n6476 ^ x200 ;
  assign n6478 = x70 ^ x32 ;
  assign n6479 = x841 ^ x96 ;
  assign n6480 = x70 & ~n6479 ;
  assign n6481 = n6480 ^ x841 ;
  assign n6482 = ~n1537 & n1782 ;
  assign n6483 = n6482 ^ x198 ;
  assign n6484 = n6483 ^ x70 ;
  assign n6485 = n6484 ^ n6478 ;
  assign n6486 = ~n6481 & n6485 ;
  assign n6487 = n6486 ^ x70 ;
  assign n6488 = n6478 & n6487 ;
  assign n6489 = ~x233 & n6488 ;
  assign n6490 = n6489 ^ n6488 ;
  assign n6491 = ~x237 & n6490 ;
  assign n6492 = n6491 ^ n6490 ;
  assign n6493 = ~x332 & ~n1323 ;
  assign n6494 = n1247 & n4210 ;
  assign n6495 = n6493 & n6494 ;
  assign n6496 = n6495 ^ n6493 ;
  assign n6497 = ~n6492 & n6496 ;
  assign n6498 = x947 ^ x587 ;
  assign n6499 = n1537 & n2655 ;
  assign n6500 = n6498 & n6499 ;
  assign n6501 = n6500 ^ n2879 ;
  assign n6502 = ~x332 & ~n6501 ;
  assign n6503 = x96 & n6483 ;
  assign n6504 = ~x237 & n6503 ;
  assign n6505 = n6504 ^ n6503 ;
  assign n6506 = ~x233 & n6501 ;
  assign n6507 = n6506 ^ n6501 ;
  assign n6508 = n6505 & n6507 ;
  assign n6509 = ~x201 & ~n6508 ;
  assign n6510 = ~n6502 & n6509 ;
  assign n6511 = ~n6497 & n6510 ;
  assign n6512 = n6511 ^ n6509 ;
  assign n6513 = n6512 ^ n6508 ;
  assign n6514 = ~x237 & n6489 ;
  assign n6515 = n6514 ^ n6489 ;
  assign n6516 = n6496 & ~n6515 ;
  assign n6517 = n6505 & n6506 ;
  assign n6518 = ~x202 & ~n6517 ;
  assign n6519 = ~n6516 & n6518 ;
  assign n6520 = ~n6502 & n6519 ;
  assign n6521 = n6520 ^ n6518 ;
  assign n6522 = n6521 ^ n6517 ;
  assign n6523 = n6496 & ~n6514 ;
  assign n6524 = n6504 & n6506 ;
  assign n6525 = ~x203 & ~n6524 ;
  assign n6526 = ~n6523 & n6525 ;
  assign n6527 = ~n6502 & n6526 ;
  assign n6528 = n6527 ^ n6525 ;
  assign n6529 = n6528 ^ n6524 ;
  assign n6531 = n2668 ^ x602 ;
  assign n6530 = n2668 ^ x907 ;
  assign n6532 = n6531 ^ n6530 ;
  assign n6535 = n1537 & n6532 ;
  assign n6536 = n6535 ^ n6530 ;
  assign n6537 = n2655 & n6536 ;
  assign n6538 = n6537 ^ n2668 ;
  assign n6539 = ~x332 & ~n6538 ;
  assign n6540 = n6505 & n6538 ;
  assign n6541 = ~x233 & n6540 ;
  assign n6542 = n6541 ^ n6540 ;
  assign n6543 = ~x204 & ~n6542 ;
  assign n6544 = ~n6539 & n6543 ;
  assign n6545 = ~n6497 & n6544 ;
  assign n6546 = n6545 ^ n6543 ;
  assign n6547 = n6546 ^ n6542 ;
  assign n6548 = ~x205 & ~n6541 ;
  assign n6549 = ~n6539 & n6548 ;
  assign n6550 = ~n6516 & n6549 ;
  assign n6551 = n6550 ^ n6548 ;
  assign n6552 = n6551 ^ n6541 ;
  assign n6553 = ~n6491 & n6496 ;
  assign n6554 = n6504 & n6538 ;
  assign n6555 = ~x233 & n6554 ;
  assign n6556 = n6555 ^ n6554 ;
  assign n6557 = ~x206 & ~n6556 ;
  assign n6558 = ~n6553 & n6557 ;
  assign n6559 = ~n6539 & n6558 ;
  assign n6560 = n6559 ^ n6557 ;
  assign n6561 = n6560 ^ n6556 ;
  assign n6569 = x623 ^ x207 ;
  assign n6566 = x710 & n5838 ;
  assign n6567 = n6566 ^ x623 ;
  assign n6568 = ~n5802 & n6567 ;
  assign n6570 = n6569 ^ n6568 ;
  assign n6571 = n5766 & ~n6570 ;
  assign n6572 = n6571 ^ x207 ;
  assign n6580 = x607 ^ x208 ;
  assign n6577 = x638 & n5838 ;
  assign n6578 = n6577 ^ x607 ;
  assign n6579 = ~n5802 & n6578 ;
  assign n6581 = n6580 ^ n6579 ;
  assign n6582 = n5766 & ~n6581 ;
  assign n6583 = n6582 ^ x208 ;
  assign n6591 = x622 ^ x209 ;
  assign n6588 = x639 & n5838 ;
  assign n6589 = n6588 ^ x622 ;
  assign n6590 = ~n5802 & n6589 ;
  assign n6592 = n6591 ^ n6590 ;
  assign n6593 = n5766 & ~n6592 ;
  assign n6594 = n6593 ^ x209 ;
  assign n6600 = x633 ^ x210 ;
  assign n6597 = x634 & x907 ;
  assign n6598 = n6597 ^ x633 ;
  assign n6599 = ~x947 & n6598 ;
  assign n6601 = n6600 ^ n6599 ;
  assign n6602 = n5766 & n6601 ;
  assign n6603 = n6602 ^ x210 ;
  assign n6609 = x606 ^ x211 ;
  assign n6606 = x643 & x907 ;
  assign n6607 = n6606 ^ x606 ;
  assign n6608 = ~x947 & n6607 ;
  assign n6610 = n6609 ^ n6608 ;
  assign n6611 = n5766 & n6610 ;
  assign n6612 = n6611 ^ x211 ;
  assign n6620 = ~x212 & ~n5766 ;
  assign n6615 = x638 & x907 ;
  assign n6616 = n6615 ^ x607 ;
  assign n6617 = ~x947 & n6616 ;
  assign n6618 = n6617 ^ x607 ;
  assign n6619 = n5943 & n6618 ;
  assign n6622 = n6620 ^ n6619 ;
  assign n6630 = ~x213 & ~n5766 ;
  assign n6625 = x639 & x907 ;
  assign n6626 = n6625 ^ x622 ;
  assign n6627 = ~x947 & n6626 ;
  assign n6628 = n6627 ^ x622 ;
  assign n6629 = n5943 & n6628 ;
  assign n6632 = n6630 ^ n6629 ;
  assign n6638 = x623 ^ x214 ;
  assign n6635 = x710 & x907 ;
  assign n6636 = n6635 ^ x623 ;
  assign n6637 = ~x947 & n6636 ;
  assign n6639 = n6638 ^ n6637 ;
  assign n6640 = n5766 & ~n6639 ;
  assign n6641 = n6640 ^ x214 ;
  assign n6649 = x642 ^ x215 ;
  assign n6646 = x681 & x907 ;
  assign n6647 = n6646 ^ x642 ;
  assign n6648 = ~x947 & n6647 ;
  assign n6650 = n6649 ^ n6648 ;
  assign n6651 = n5766 & n6650 ;
  assign n6652 = n6651 ^ x215 ;
  assign n6660 = x614 ^ x216 ;
  assign n6657 = x662 & x907 ;
  assign n6658 = n6657 ^ x614 ;
  assign n6659 = ~x947 & n6658 ;
  assign n6661 = n6660 ^ n6659 ;
  assign n6662 = n5766 & n6661 ;
  assign n6663 = n6662 ^ x216 ;
  assign n6671 = x612 ^ x217 ;
  assign n6668 = ~x695 & n5838 ;
  assign n6669 = n6668 ^ x612 ;
  assign n6670 = ~n5802 & n6669 ;
  assign n6672 = n6671 ^ n6670 ;
  assign n6673 = n5766 & ~n6672 ;
  assign n6674 = n6673 ^ x217 ;
  assign n6675 = ~x218 & ~n6555 ;
  assign n6676 = ~n6539 & n6675 ;
  assign n6677 = ~n6523 & n6676 ;
  assign n6678 = n6677 ^ n6675 ;
  assign n6679 = n6678 ^ n6555 ;
  assign n6687 = x219 & ~n5766 ;
  assign n6682 = x637 & x907 ;
  assign n6683 = n6682 ^ x617 ;
  assign n6684 = ~x947 & n6683 ;
  assign n6685 = n6684 ^ x617 ;
  assign n6686 = n5943 & n6685 ;
  assign n6689 = n6687 ^ n6686 ;
  assign n6690 = n6504 & n6507 ;
  assign n6691 = ~x220 & ~n6690 ;
  assign n6692 = ~n6553 & n6691 ;
  assign n6693 = ~n6502 & n6692 ;
  assign n6694 = n6693 ^ n6691 ;
  assign n6695 = n6694 ^ n6690 ;
  assign n6703 = x616 ^ x221 ;
  assign n6700 = x661 & x907 ;
  assign n6701 = n6700 ^ x616 ;
  assign n6702 = ~x947 & n6701 ;
  assign n6704 = n6703 ^ n6702 ;
  assign n6705 = n5766 & n6704 ;
  assign n6706 = n6705 ^ x221 ;
  assign n6712 = x616 ^ x222 ;
  assign n6709 = x661 & n5838 ;
  assign n6710 = n6709 ^ x616 ;
  assign n6711 = ~n5802 & n6710 ;
  assign n6713 = n6712 ^ n6711 ;
  assign n6714 = n5766 & n6713 ;
  assign n6715 = n6714 ^ x222 ;
  assign n6721 = x642 ^ x223 ;
  assign n6718 = x681 & n5838 ;
  assign n6719 = n6718 ^ x642 ;
  assign n6720 = ~n5802 & n6719 ;
  assign n6722 = n6721 ^ n6720 ;
  assign n6723 = n5766 & n6722 ;
  assign n6724 = n6723 ^ x223 ;
  assign n6730 = x614 ^ x224 ;
  assign n6727 = x662 & n5838 ;
  assign n6728 = n6727 ^ x614 ;
  assign n6729 = ~n5802 & n6728 ;
  assign n6731 = n6730 ^ n6729 ;
  assign n6732 = n5766 & n6731 ;
  assign n6733 = n6732 ^ x224 ;
  assign n6754 = n1556 & n1880 ;
  assign n6734 = ~n1788 & n1919 ;
  assign n6735 = x70 & n6734 ;
  assign n6736 = x332 & n6735 ;
  assign n6737 = n6736 ^ n6734 ;
  assign n6738 = n6737 ^ n1919 ;
  assign n6739 = ~x55 & ~x137 ;
  assign n6740 = ~n1341 & n6739 ;
  assign n6749 = n1798 & n5065 ;
  assign n6750 = n6740 & n6749 ;
  assign n6751 = n6750 ^ n6740 ;
  assign n6752 = n6751 ^ n1341 ;
  assign n6753 = ~n6738 & n6752 ;
  assign n6756 = n6754 ^ n6753 ;
  assign n6759 = ~n1292 & n1338 ;
  assign n6757 = x479 & n4819 ;
  assign n6758 = n6757 ^ n1304 ;
  assign n6761 = n6759 ^ n6758 ;
  assign n6762 = n1919 & ~n6761 ;
  assign n6763 = n2740 & n6762 ;
  assign n6764 = n6763 ^ n6761 ;
  assign n6765 = n6764 ^ x231 ;
  assign n6766 = ~x228 & n6765 ;
  assign n6767 = n6766 ^ x231 ;
  assign n6768 = n1564 & n1816 ;
  assign n6769 = ~x58 & n6768 ;
  assign n6770 = n6769 ^ x72 ;
  assign n6771 = ~x72 & ~n6770 ;
  assign n6772 = n4138 & n6771 ;
  assign n6773 = n1919 & n6772 ;
  assign n6781 = x1093 & n6773 ;
  assign n6782 = n3927 & n6781 ;
  assign n6783 = n6782 ^ n3927 ;
  assign n6774 = n6773 ^ n1919 ;
  assign n6775 = n6774 ^ n3927 ;
  assign n6784 = n6783 ^ n6775 ;
  assign n6785 = ~n4377 & ~n6784 ;
  assign n6786 = x36 & n1851 ;
  assign n6787 = ~n6785 & n6786 ;
  assign n6788 = n6787 ^ n6785 ;
  assign n6795 = x1091 & n4756 ;
  assign n6789 = n1280 & n1290 ;
  assign n6790 = n1863 ^ n1846 ;
  assign n6791 = n1860 & n6790 ;
  assign n6792 = n6789 & n6791 ;
  assign n6793 = ~x228 & ~n6792 ;
  assign n6794 = ~x39 & ~n6793 ;
  assign n6797 = n6795 ^ n6794 ;
  assign n6798 = ~x47 & n1245 ;
  assign n6799 = ~n2608 & ~n3537 ;
  assign n6800 = n6798 & n6799 ;
  assign n6801 = ~n5765 & ~n6800 ;
  assign n6842 = n4321 ^ n3886 ;
  assign n6803 = n4321 ^ n1341 ;
  assign n6843 = n6842 ^ n6803 ;
  assign n6808 = x102 ^ x65 ;
  assign n6809 = ~x64 & n3539 ;
  assign n6810 = n1638 & n6809 ;
  assign n6811 = n6808 & n6810 ;
  assign n6846 = n6843 ^ n6811 ;
  assign n6844 = n6843 ^ n2761 ;
  assign n6845 = n6844 ^ n6803 ;
  assign n6864 = n6846 ^ n6845 ;
  assign n6865 = n6864 ^ n6842 ;
  assign n6866 = n6865 ^ n4321 ;
  assign n6847 = n6846 ^ n6803 ;
  assign n6848 = n6847 ^ n6845 ;
  assign n6830 = n6865 ^ n1341 ;
  assign n6816 = n6864 ^ n6843 ;
  assign n6832 = n6846 ^ n6816 ;
  assign n6831 = ~n6830 & n6832 ;
  assign n6838 = n6831 ^ n4321 ;
  assign n6839 = n6848 ^ n6838 ;
  assign n6860 = n6839 ^ n3886 ;
  assign n6861 = n6866 ^ n6860 ;
  assign n6862 = n6861 ^ n6848 ;
  assign n6869 = n6862 ^ n3886 ;
  assign n6870 = n6869 ^ n1341 ;
  assign n6871 = n6870 ^ n6866 ;
  assign n6872 = x209 & n1537 ;
  assign n6873 = n6872 ^ n1537 ;
  assign n6897 = x1155 & ~n4362 ;
  assign n6896 = x1153 & n4074 ;
  assign n6898 = n6897 ^ n6896 ;
  assign n6895 = x1154 & n4092 ;
  assign n6899 = n6898 ^ n6895 ;
  assign n6900 = x208 & n6899 ;
  assign n6874 = x1156 ^ x1155 ;
  assign n6875 = x200 & n6874 ;
  assign n6876 = n6875 ^ x1155 ;
  assign n6886 = n6876 ^ n6874 ;
  assign n6887 = ~x199 & n6886 ;
  assign n6885 = x1154 & n4074 ;
  assign n6888 = n6887 ^ n6885 ;
  assign n6881 = ~x200 & x1157 ;
  assign n6882 = n6881 ^ n6876 ;
  assign n6883 = ~n4091 & n6882 ;
  assign n6884 = n6883 ^ n6876 ;
  assign n6889 = n6888 ^ n6884 ;
  assign n6890 = x207 & n6889 ;
  assign n6891 = n6890 ^ n6888 ;
  assign n6901 = n6900 ^ n6891 ;
  assign n6923 = n4075 ^ x208 ;
  assign n7194 = n6923 ^ n4076 ;
  assign n6902 = n6901 & ~n7194 ;
  assign n6903 = n6902 ^ n6891 ;
  assign n6904 = n6873 & n6903 ;
  assign n6905 = n6904 ^ n6873 ;
  assign n6960 = x1155 ^ x1154 ;
  assign n6963 = ~x214 & n6960 ;
  assign n6964 = n6963 ^ x1154 ;
  assign n6965 = ~x219 & n6964 ;
  assign n6940 = x1156 ^ x1154 ;
  assign n6941 = ~x219 & n6940 ;
  assign n6942 = n6941 ^ x1154 ;
  assign n6937 = x1155 ^ x1153 ;
  assign n6938 = ~x219 & n6937 ;
  assign n6939 = n6938 ^ x1153 ;
  assign n6943 = n6942 ^ n6939 ;
  assign n6944 = x214 & n6943 ;
  assign n6945 = n6944 ^ n6942 ;
  assign n6966 = n6965 ^ n6945 ;
  assign n6967 = x211 & n6966 ;
  assign n6946 = x214 ^ x212 ;
  assign n6947 = ~x219 & n6946 ;
  assign n6948 = x211 & n6947 ;
  assign n6955 = n6948 ^ n6947 ;
  assign n6956 = x1144 & n6955 ;
  assign n6952 = ~n4071 & n4084 ;
  assign n6951 = ~n4073 & n4083 ;
  assign n6953 = n6952 ^ n6951 ;
  assign n6954 = x1142 & n6953 ;
  assign n6957 = n6956 ^ n6954 ;
  assign n6949 = n6948 ^ n4249 ;
  assign n6950 = x1143 & n6949 ;
  assign n6958 = n6957 ^ n6950 ;
  assign n6959 = n6958 ^ n6945 ;
  assign n6968 = n6967 ^ n6959 ;
  assign n6979 = n6968 ^ n6958 ;
  assign n6974 = ~x219 & x1156 ;
  assign n6969 = x1157 ^ x1155 ;
  assign n6970 = ~x219 & n6969 ;
  assign n6971 = n6970 ^ x1155 ;
  assign n6975 = n6974 ^ n6971 ;
  assign n6976 = x211 & n6975 ;
  assign n6977 = n6976 ^ n6971 ;
  assign n6978 = x214 & n6977 ;
  assign n6980 = n6979 ^ n6978 ;
  assign n6981 = ~x212 & n6980 ;
  assign n6982 = n6981 ^ n6968 ;
  assign n6983 = ~x213 & n6982 ;
  assign n6984 = n6983 ^ n6958 ;
  assign n6985 = ~n1537 & ~n6984 ;
  assign n6906 = x1142 & ~n4245 ;
  assign n6907 = n7194 ^ x200 ;
  assign n6912 = x1144 & n7194 ;
  assign n6913 = n6912 ^ x1143 ;
  assign n6914 = ~n6907 & n6913 ;
  assign n6919 = ~x208 & n6914 ;
  assign n6920 = n6919 ^ x1144 ;
  assign n6921 = n6920 & ~n7194 ;
  assign n6915 = n6914 ^ x1144 ;
  assign n6922 = n6921 ^ n6915 ;
  assign n6933 = n4362 & ~n6922 ;
  assign n6934 = n6906 & n6933 ;
  assign n6924 = ~x200 & n6923 ;
  assign n6925 = n6924 ^ n6922 ;
  assign n6928 = ~x1142 & ~n6925 ;
  assign n6929 = n6928 ^ n6924 ;
  assign n6930 = x199 & ~n6929 ;
  assign n6931 = n6930 ^ n6922 ;
  assign n6935 = n6934 ^ n6931 ;
  assign n6936 = n6872 & ~n6935 ;
  assign n6986 = n6985 ^ n6936 ;
  assign n6987 = ~n6905 & ~n6986 ;
  assign n6988 = n6987 ^ x233 ;
  assign n6989 = x230 & ~n6988 ;
  assign n6990 = n6989 ^ x233 ;
  assign n7011 = n6923 ^ n4071 ;
  assign n7012 = n1537 & ~n7011 ;
  assign n7013 = n7012 ^ n4071 ;
  assign n7023 = n4100 & ~n4252 ;
  assign n7024 = ~n7013 & n7023 ;
  assign n7025 = x1152 & n7024 ;
  assign n7014 = ~n4100 & ~n7013 ;
  assign n7015 = x1154 ^ x1153 ;
  assign n7020 = n4252 & n7015 ;
  assign n7021 = n7020 ^ x1153 ;
  assign n7022 = n7014 & n7021 ;
  assign n7027 = n7025 ^ n7022 ;
  assign n7039 = n7027 ^ x234 ;
  assign n6991 = x213 & ~n1537 ;
  assign n6993 = x1156 & n6955 ;
  assign n6994 = n6991 & n6993 ;
  assign n6995 = n6994 ^ x1155 ;
  assign n6996 = n6994 ^ n6991 ;
  assign n7006 = n6949 & n6996 ;
  assign n7007 = n6995 & n7006 ;
  assign n7008 = n7007 ^ n6996 ;
  assign n6999 = x208 & n6897 ;
  assign n7000 = n6999 ^ n6887 ;
  assign n7001 = n7000 & ~n7194 ;
  assign n7002 = n7001 ^ n6887 ;
  assign n7003 = n6872 & n7002 ;
  assign n7004 = n7003 ^ n6872 ;
  assign n7009 = n7008 ^ n7004 ;
  assign n7040 = n7039 ^ n7009 ;
  assign n6992 = n6991 ^ n6872 ;
  assign n7041 = n7040 ^ n6992 ;
  assign n7033 = x1154 & n7024 ;
  assign n7028 = n7027 ^ n6992 ;
  assign n7034 = n7033 ^ n7028 ;
  assign n7035 = n7009 & ~n7034 ;
  assign n7042 = n7041 ^ n7035 ;
  assign n7010 = n7009 ^ n6992 ;
  assign n7036 = n7027 ^ n7009 ;
  assign n7037 = ~n7035 & n7036 ;
  assign n7038 = n7010 & n7037 ;
  assign n7043 = n7042 ^ n7038 ;
  assign n7044 = x230 & n7043 ;
  assign n7045 = n7044 ^ x234 ;
  assign n7046 = n1537 & n4076 ;
  assign n7049 = ~x200 & n7015 ;
  assign n7050 = n7049 ^ x1153 ;
  assign n7051 = ~x199 & n7050 ;
  assign n7052 = n7051 ^ n6887 ;
  assign n7055 = ~x209 & n7052 ;
  assign n7056 = n7055 ^ n6887 ;
  assign n7057 = n7046 & n7056 ;
  assign n7058 = n7057 ^ n1537 ;
  assign n7059 = n7058 & n7194 ;
  assign n7060 = n6899 ^ n6884 ;
  assign n7063 = x209 & n7060 ;
  assign n7064 = n7063 ^ n6899 ;
  assign n7065 = n7059 & n7064 ;
  assign n7066 = n7065 ^ n7058 ;
  assign n7067 = ~n1537 & n6951 ;
  assign n7070 = ~x213 & n6937 ;
  assign n7071 = n7070 ^ x1155 ;
  assign n7072 = n7067 & n7071 ;
  assign n7073 = n7072 ^ n1537 ;
  assign n7074 = ~x211 & n6946 ;
  assign n7075 = n6971 ^ n6939 ;
  assign n7078 = x213 & n7075 ;
  assign n7079 = n7078 ^ n6939 ;
  assign n7080 = n7074 & n7079 ;
  assign n7081 = ~n7073 & ~n7080 ;
  assign n7082 = n6949 & n7081 ;
  assign n7085 = ~x213 & n6940 ;
  assign n7086 = n7085 ^ x1156 ;
  assign n7087 = n7082 & n7086 ;
  assign n7088 = n7087 ^ n7081 ;
  assign n7089 = ~n7066 & ~n7088 ;
  assign n7090 = n7089 ^ x235 ;
  assign n7091 = x230 & n7090 ;
  assign n7092 = n7091 ^ x235 ;
  assign n7173 = x208 & n6888 ;
  assign n7160 = ~x200 & x1158 ;
  assign n7113 = x1157 ^ x1156 ;
  assign n7154 = x200 & n7113 ;
  assign n7155 = n7154 ^ x1156 ;
  assign n7161 = n7160 ^ n7155 ;
  assign n7162 = ~n4091 & n7161 ;
  assign n7163 = n7162 ^ n7155 ;
  assign n7164 = n7163 ^ n6884 ;
  assign n7165 = ~x208 & n7164 ;
  assign n7166 = n7165 ^ n6884 ;
  assign n7174 = n7173 ^ n7166 ;
  assign n7175 = n7174 & ~n7194 ;
  assign n7149 = n7194 ^ n6924 ;
  assign n7150 = ~x199 & x1144 ;
  assign n7151 = n7149 & n7150 ;
  assign n7139 = ~x199 & n4076 ;
  assign n7140 = n7139 ^ n6924 ;
  assign n7141 = x1145 ^ x1143 ;
  assign n7143 = n4245 & n7141 ;
  assign n7144 = n7143 ^ x1145 ;
  assign n7145 = n7144 ^ n7141 ;
  assign n7146 = ~n7140 & n7145 ;
  assign n7147 = n7146 ^ n7143 ;
  assign n7148 = n7147 ^ x1143 ;
  assign n7152 = n7151 ^ n7148 ;
  assign n7167 = n7166 ^ n7152 ;
  assign n7176 = n7175 ^ n7167 ;
  assign n7177 = ~x209 & n7176 ;
  assign n7114 = ~x219 & n7113 ;
  assign n7106 = n6971 ^ n6942 ;
  assign n7107 = ~x214 & n7106 ;
  assign n7108 = n7107 ^ n6942 ;
  assign n7103 = ~x214 & n6874 ;
  assign n7104 = n7103 ^ x1155 ;
  assign n7105 = ~x219 & n7104 ;
  assign n7109 = n7108 ^ n7105 ;
  assign n7110 = x211 & n7109 ;
  assign n7111 = n7110 ^ n7108 ;
  assign n7095 = x1158 ^ x1157 ;
  assign n7096 = n7095 ^ x1156 ;
  assign n7097 = ~x219 & n7096 ;
  assign n7098 = n7097 ^ x1156 ;
  assign n7099 = ~n4082 & n7098 ;
  assign n7100 = n7099 ^ x1156 ;
  assign n7112 = n7111 ^ n7100 ;
  assign n7115 = n7114 ^ n7112 ;
  assign n7223 = n7115 ^ n7111 ;
  assign n7126 = ~x214 & n7223 ;
  assign n7127 = n7126 ^ n7115 ;
  assign n7128 = ~x212 & n7127 ;
  assign n7121 = x1143 & n6953 ;
  assign n7119 = x1145 & n6955 ;
  assign n7118 = x1144 & n6949 ;
  assign n7120 = n7119 ^ n7118 ;
  assign n7122 = n7121 ^ n7120 ;
  assign n7123 = n7122 ^ n7111 ;
  assign n7129 = n7128 ^ n7123 ;
  assign n7130 = ~x213 & n7129 ;
  assign n7131 = n7130 ^ n7122 ;
  assign n7153 = n7152 ^ n7131 ;
  assign n7178 = n7177 ^ n7153 ;
  assign n7179 = n1537 & n7178 ;
  assign n7132 = n7131 ^ x237 ;
  assign n7180 = n7179 ^ n7132 ;
  assign n7181 = x230 & ~n7180 ;
  assign n7182 = n7181 ^ x237 ;
  assign n7202 = x1154 & n6949 ;
  assign n7201 = x1155 & n6955 ;
  assign n7203 = n7202 ^ n7201 ;
  assign n7200 = x1153 & n6953 ;
  assign n7204 = n7203 ^ n7200 ;
  assign n7205 = n6991 & ~n7204 ;
  assign n7209 = n7205 ^ x238 ;
  assign n7191 = n6872 & n6899 ;
  assign n7196 = n4076 & ~n6896 ;
  assign n7197 = n7196 ^ n6923 ;
  assign n7198 = n7191 & n7197 ;
  assign n7199 = n7198 ^ n6872 ;
  assign n7210 = n7209 ^ n7199 ;
  assign n7207 = n4076 & n7199 ;
  assign n7208 = n7051 & n7207 ;
  assign n7211 = n7210 ^ n7208 ;
  assign n7187 = x1151 & n7024 ;
  assign n7183 = x1153 ^ x1152 ;
  assign n7184 = ~n4252 & n7183 ;
  assign n7185 = n7184 ^ x1153 ;
  assign n7186 = n7014 & n7185 ;
  assign n7189 = n7187 ^ n7186 ;
  assign n7190 = ~n6992 & ~n7189 ;
  assign n7212 = n7211 ^ n7190 ;
  assign n7213 = x230 & ~n7212 ;
  assign n7214 = n7213 ^ x238 ;
  assign n7215 = n1537 & n4075 ;
  assign n7216 = n7163 ^ n6888 ;
  assign n7219 = x209 & n7216 ;
  assign n7220 = n7219 ^ n6888 ;
  assign n7221 = n7215 & n7220 ;
  assign n7222 = ~n1537 & ~n4072 ;
  assign n7227 = x213 & n7115 ;
  assign n7228 = n7227 ^ n7111 ;
  assign n7229 = n7222 & n7228 ;
  assign n7230 = ~n7221 & ~n7229 ;
  assign n7231 = n7230 ^ x239 ;
  assign n7232 = x230 & ~n7231 ;
  assign n7233 = n7232 ^ x239 ;
  assign n7252 = x1147 & n7024 ;
  assign n7246 = x1149 ^ x1148 ;
  assign n7249 = ~n4252 & n7246 ;
  assign n7250 = n7249 ^ x1149 ;
  assign n7251 = n7014 & n7250 ;
  assign n7254 = n7252 ^ n7251 ;
  assign n7255 = n7254 ^ x240 ;
  assign n7240 = x1145 & n7024 ;
  assign n7234 = x1147 ^ x1146 ;
  assign n7237 = ~n4252 & n7234 ;
  assign n7238 = n7237 ^ x1147 ;
  assign n7239 = n7014 & n7238 ;
  assign n7242 = n7240 ^ n7239 ;
  assign n7243 = n7242 ^ x240 ;
  assign n7256 = n7255 ^ n7243 ;
  assign n7257 = n6992 & n7256 ;
  assign n7258 = n7257 ^ n7243 ;
  assign n7259 = x230 & n7258 ;
  assign n7260 = n7259 ^ x240 ;
  assign n7270 = x1149 & n7024 ;
  assign n7264 = x1151 ^ x1150 ;
  assign n7267 = ~n4252 & n7264 ;
  assign n7268 = n7267 ^ x1151 ;
  assign n7269 = n7014 & n7268 ;
  assign n7272 = n7270 ^ n7269 ;
  assign n7273 = n7272 ^ x241 ;
  assign n7261 = n7189 ^ x241 ;
  assign n7274 = n7273 ^ n7261 ;
  assign n7275 = ~n6992 & n7274 ;
  assign n7276 = n7275 ^ n7261 ;
  assign n7277 = x230 & n7276 ;
  assign n7278 = n7277 ^ x241 ;
  assign n7291 = n6873 & ~n6935 ;
  assign n7287 = x1144 & n7024 ;
  assign n7281 = x1146 ^ x1145 ;
  assign n7284 = ~n4252 & n7281 ;
  assign n7285 = n7284 ^ x1146 ;
  assign n7286 = n7014 & n7285 ;
  assign n7289 = n7287 ^ n7286 ;
  assign n7290 = n6992 & ~n7289 ;
  assign n7292 = n7291 ^ n7290 ;
  assign n7293 = n7292 ^ x242 ;
  assign n7279 = n6991 ^ n1537 ;
  assign n7280 = ~n6958 & ~n7279 ;
  assign n7294 = n7293 ^ n7280 ;
  assign n7295 = x230 & ~n7294 ;
  assign n7296 = n7295 ^ x242 ;
  assign n7297 = ~x230 & ~x1091 ;
  assign n7322 = n4099 ^ n4095 ;
  assign n7323 = x1155 & n7322 ;
  assign n7318 = n4084 ^ n4074 ;
  assign n7319 = n1537 & n7318 ;
  assign n7320 = n7319 ^ n4084 ;
  assign n7321 = x1157 & n7320 ;
  assign n7324 = n7323 ^ n7321 ;
  assign n7299 = ~x83 & ~x85 ;
  assign n7300 = x314 & n7299 ;
  assign n7302 = x81 & ~n4099 ;
  assign n7303 = n7300 & n7302 ;
  assign n7301 = n7300 ^ x314 ;
  assign n7304 = n7303 ^ n7301 ;
  assign n7305 = x802 & n7304 ;
  assign n7306 = x276 & n7305 ;
  assign n7307 = x271 & n7306 ;
  assign n7308 = x273 & n7307 ;
  assign n7309 = x283 & n7308 ;
  assign n7310 = x272 & n7309 ;
  assign n7311 = x275 & n7310 ;
  assign n7312 = x268 & n7311 ;
  assign n7313 = x253 & n7312 ;
  assign n7314 = x254 & n7313 ;
  assign n7315 = x267 & n7314 ;
  assign n7316 = ~x263 & n7315 ;
  assign n7317 = n7316 ^ x243 ;
  assign n7325 = n7324 ^ n7317 ;
  assign n7298 = x1156 & ~n4095 ;
  assign n7326 = n7325 ^ n7298 ;
  assign n7327 = ~n7297 & ~n7326 ;
  assign n7328 = n7327 ^ n7317 ;
  assign n7331 = ~n7122 & ~n7279 ;
  assign n7330 = n6992 & ~n7242 ;
  assign n7332 = n7331 ^ n7330 ;
  assign n7333 = n7332 ^ x244 ;
  assign n7329 = n6873 & ~n7152 ;
  assign n7334 = n7333 ^ n7329 ;
  assign n7335 = x230 & ~n7334 ;
  assign n7336 = n7335 ^ x244 ;
  assign n7346 = x1146 & n7024 ;
  assign n7340 = x1148 ^ x1147 ;
  assign n7343 = ~n4252 & n7340 ;
  assign n7344 = n7343 ^ x1148 ;
  assign n7345 = n7014 & n7344 ;
  assign n7348 = n7346 ^ n7345 ;
  assign n7349 = n7348 ^ x245 ;
  assign n7337 = n7289 ^ x245 ;
  assign n7350 = n7349 ^ n7337 ;
  assign n7351 = n6992 & n7350 ;
  assign n7352 = n7351 ^ n7337 ;
  assign n7353 = x230 & n7352 ;
  assign n7354 = n7353 ^ x245 ;
  assign n7364 = x1148 & n7024 ;
  assign n7358 = x1150 ^ x1149 ;
  assign n7361 = ~n4252 & n7358 ;
  assign n7362 = n7361 ^ x1150 ;
  assign n7363 = n7014 & n7362 ;
  assign n7366 = n7364 ^ n7363 ;
  assign n7367 = n7366 ^ x246 ;
  assign n7355 = n7348 ^ x246 ;
  assign n7368 = n7367 ^ n7355 ;
  assign n7369 = n6992 & n7368 ;
  assign n7370 = n7369 ^ n7355 ;
  assign n7371 = x230 & n7370 ;
  assign n7372 = n7371 ^ x246 ;
  assign n7376 = n7272 ^ x247 ;
  assign n7373 = n7254 ^ x247 ;
  assign n7377 = n7376 ^ n7373 ;
  assign n7378 = n6992 & n7377 ;
  assign n7379 = n7378 ^ n7373 ;
  assign n7380 = x230 & n7379 ;
  assign n7381 = n7380 ^ x247 ;
  assign n7391 = x1150 & n7024 ;
  assign n7385 = x1152 ^ x1151 ;
  assign n7388 = ~n4252 & n7385 ;
  assign n7389 = n7388 ^ x1152 ;
  assign n7390 = n7014 & n7389 ;
  assign n7393 = n7391 ^ n7390 ;
  assign n7394 = n7393 ^ x248 ;
  assign n7382 = n7366 ^ x248 ;
  assign n7395 = n7394 ^ n7382 ;
  assign n7396 = n6992 & n7395 ;
  assign n7397 = n7396 ^ n7382 ;
  assign n7398 = x230 & n7397 ;
  assign n7399 = n7398 ^ x248 ;
  assign n7403 = n7393 ^ x249 ;
  assign n7400 = n7027 ^ x249 ;
  assign n7404 = n7403 ^ n7400 ;
  assign n7405 = ~n6992 & n7404 ;
  assign n7406 = n7405 ^ n7400 ;
  assign n7407 = x230 & n7406 ;
  assign n7408 = n7407 ^ x249 ;
  assign n7409 = ~x250 & ~n4218 ;
  assign n7410 = ~n5065 & n7409 ;
  assign n7411 = n7410 ^ x250 ;
  assign n7412 = x1053 ^ x1039 ;
  assign n7413 = ~x200 & n7412 ;
  assign n7414 = n7413 ^ x1039 ;
  assign n7415 = n7414 ^ x251 ;
  assign n7416 = x897 ^ x476 ;
  assign n7417 = ~x200 & ~n7416 ;
  assign n7418 = n7417 ^ x476 ;
  assign n7419 = ~x199 & ~n7418 ;
  assign n7420 = n7415 & n7419 ;
  assign n7421 = n7420 ^ x251 ;
  assign n7422 = n2704 & ~n2707 ;
  assign n7423 = n2966 & n7422 ;
  assign n7424 = x252 & x1092 ;
  assign n7425 = ~n7423 & n7424 ;
  assign n7427 = x1093 & ~n3209 ;
  assign n7428 = n7425 & n7427 ;
  assign n7426 = n7425 ^ n7423 ;
  assign n7429 = n7428 ^ n7426 ;
  assign n7433 = x1151 & n7322 ;
  assign n7432 = x1153 & n7320 ;
  assign n7434 = n7433 ^ n7432 ;
  assign n7431 = n7312 ^ x253 ;
  assign n7435 = n7434 ^ n7431 ;
  assign n7430 = x1152 & ~n4095 ;
  assign n7436 = n7435 ^ n7430 ;
  assign n7437 = ~n7297 & n7436 ;
  assign n7438 = n7437 ^ n7431 ;
  assign n7442 = x1154 & n7320 ;
  assign n7441 = x1152 & n7322 ;
  assign n7443 = n7442 ^ n7441 ;
  assign n7440 = n7313 ^ x254 ;
  assign n7444 = n7443 ^ n7440 ;
  assign n7439 = x1153 & ~n4095 ;
  assign n7445 = n7444 ^ n7439 ;
  assign n7446 = ~n7297 & n7445 ;
  assign n7447 = n7446 ^ n7440 ;
  assign n7448 = x1049 ^ x1036 ;
  assign n7449 = ~x200 & n7448 ;
  assign n7450 = n7449 ^ x1036 ;
  assign n7451 = n7450 ^ x255 ;
  assign n7452 = n7419 & n7451 ;
  assign n7453 = n7452 ^ x255 ;
  assign n7454 = x1070 ^ x1048 ;
  assign n7455 = x200 & n7454 ;
  assign n7456 = n7455 ^ x1048 ;
  assign n7457 = n7456 ^ x256 ;
  assign n7458 = n7419 & n7457 ;
  assign n7459 = n7458 ^ x256 ;
  assign n7460 = x1084 ^ x1065 ;
  assign n7461 = ~x200 & n7460 ;
  assign n7462 = n7461 ^ x1065 ;
  assign n7463 = n7462 ^ x257 ;
  assign n7464 = n7419 & n7463 ;
  assign n7465 = n7464 ^ x257 ;
  assign n7466 = x1072 ^ x1062 ;
  assign n7467 = ~x200 & n7466 ;
  assign n7468 = n7467 ^ x1062 ;
  assign n7469 = n7468 ^ x258 ;
  assign n7470 = n7419 & n7469 ;
  assign n7471 = n7470 ^ x258 ;
  assign n7472 = x1069 ^ x1059 ;
  assign n7473 = x200 & n7472 ;
  assign n7474 = n7473 ^ x1059 ;
  assign n7475 = n7474 ^ x259 ;
  assign n7476 = n7419 & n7475 ;
  assign n7477 = n7476 ^ x259 ;
  assign n7478 = x1067 ^ x1044 ;
  assign n7479 = x200 & n7478 ;
  assign n7480 = n7479 ^ x1044 ;
  assign n7481 = n7480 ^ x260 ;
  assign n7482 = n7419 & n7481 ;
  assign n7483 = n7482 ^ x260 ;
  assign n7484 = x1040 ^ x1037 ;
  assign n7485 = x200 & n7484 ;
  assign n7486 = n7485 ^ x1037 ;
  assign n7487 = n7486 ^ x261 ;
  assign n7488 = n7419 & n7487 ;
  assign n7489 = n7488 ^ x261 ;
  assign n7490 = x1093 ^ x123 ;
  assign n7491 = ~x228 & ~n7490 ;
  assign n7492 = n7491 ^ x123 ;
  assign n7497 = x1142 & n7014 ;
  assign n7498 = n7497 ^ x262 ;
  assign n7499 = ~n7492 & ~n7498 ;
  assign n7500 = n7499 ^ x262 ;
  assign n7504 = x1154 & n7322 ;
  assign n7503 = x1156 & n7320 ;
  assign n7505 = n7504 ^ n7503 ;
  assign n7502 = n7315 ^ x263 ;
  assign n7506 = n7505 ^ n7502 ;
  assign n7501 = x1155 & ~n4095 ;
  assign n7507 = n7506 ^ n7501 ;
  assign n7508 = ~n7297 & ~n7507 ;
  assign n7509 = n7508 ^ n7502 ;
  assign n7515 = x1143 & n7320 ;
  assign n7514 = x1141 & n7322 ;
  assign n7516 = n7515 ^ n7514 ;
  assign n7511 = x796 ^ x264 ;
  assign n7512 = n7304 & ~n7511 ;
  assign n7513 = n7512 ^ x264 ;
  assign n7517 = n7516 ^ n7513 ;
  assign n7510 = x1142 & ~n4095 ;
  assign n7518 = n7517 ^ n7510 ;
  assign n7519 = ~n7297 & ~n7518 ;
  assign n7520 = n7519 ^ n7513 ;
  assign n7526 = x1144 & n7320 ;
  assign n7525 = x1142 & n7322 ;
  assign n7527 = n7526 ^ n7525 ;
  assign n7522 = x819 ^ x265 ;
  assign n7523 = n7304 & ~n7522 ;
  assign n7524 = n7523 ^ x265 ;
  assign n7528 = n7527 ^ n7524 ;
  assign n7521 = x1143 & ~n4095 ;
  assign n7529 = n7528 ^ n7521 ;
  assign n7530 = ~n7297 & ~n7529 ;
  assign n7531 = n7530 ^ n7524 ;
  assign n7537 = x1136 & n7320 ;
  assign n7536 = x1134 & n7322 ;
  assign n7538 = n7537 ^ n7536 ;
  assign n7533 = x948 ^ x266 ;
  assign n7534 = n7304 & n7533 ;
  assign n7535 = n7534 ^ x266 ;
  assign n7539 = n7538 ^ n7535 ;
  assign n7532 = x1135 & ~n4095 ;
  assign n7540 = n7539 ^ n7532 ;
  assign n7541 = ~n7297 & n7540 ;
  assign n7542 = n7541 ^ n7535 ;
  assign n7546 = x1155 & n7320 ;
  assign n7545 = x1153 & n7322 ;
  assign n7547 = n7546 ^ n7545 ;
  assign n7544 = n7314 ^ x267 ;
  assign n7548 = n7547 ^ n7544 ;
  assign n7543 = x1154 & ~n4095 ;
  assign n7549 = n7548 ^ n7543 ;
  assign n7550 = ~n7297 & n7549 ;
  assign n7551 = n7550 ^ n7544 ;
  assign n7555 = x1150 & n7322 ;
  assign n7554 = x1152 & n7320 ;
  assign n7556 = n7555 ^ n7554 ;
  assign n7553 = n7311 ^ x268 ;
  assign n7557 = n7556 ^ n7553 ;
  assign n7552 = x1151 & ~n4095 ;
  assign n7558 = n7557 ^ n7552 ;
  assign n7559 = ~n7297 & n7558 ;
  assign n7560 = n7559 ^ n7553 ;
  assign n7566 = x1138 & n7320 ;
  assign n7565 = x1136 & n7322 ;
  assign n7567 = n7566 ^ n7565 ;
  assign n7562 = x817 ^ x269 ;
  assign n7563 = n7304 & ~n7562 ;
  assign n7564 = n7563 ^ x269 ;
  assign n7568 = n7567 ^ n7564 ;
  assign n7561 = x1137 & ~n4095 ;
  assign n7569 = n7568 ^ n7561 ;
  assign n7570 = ~n7297 & ~n7569 ;
  assign n7571 = n7570 ^ n7564 ;
  assign n7577 = x1141 & n7320 ;
  assign n7576 = x1139 & n7322 ;
  assign n7578 = n7577 ^ n7576 ;
  assign n7573 = x805 ^ x270 ;
  assign n7574 = n7304 & ~n7573 ;
  assign n7575 = n7574 ^ x270 ;
  assign n7579 = n7578 ^ n7575 ;
  assign n7572 = x1140 & ~n4095 ;
  assign n7580 = n7579 ^ n7572 ;
  assign n7581 = ~n7297 & ~n7580 ;
  assign n7582 = n7581 ^ n7575 ;
  assign n7586 = x1147 & n7320 ;
  assign n7585 = x1145 & n7322 ;
  assign n7587 = n7586 ^ n7585 ;
  assign n7584 = n7306 ^ x271 ;
  assign n7588 = n7587 ^ n7584 ;
  assign n7583 = x1146 & ~n4095 ;
  assign n7589 = n7588 ^ n7583 ;
  assign n7590 = ~n7297 & n7589 ;
  assign n7591 = n7590 ^ n7584 ;
  assign n7595 = x1148 & n7322 ;
  assign n7594 = x1150 & n7320 ;
  assign n7596 = n7595 ^ n7594 ;
  assign n7593 = n7309 ^ x272 ;
  assign n7597 = n7596 ^ n7593 ;
  assign n7592 = x1149 & ~n4095 ;
  assign n7598 = n7597 ^ n7592 ;
  assign n7599 = ~n7297 & n7598 ;
  assign n7600 = n7599 ^ n7593 ;
  assign n7604 = x1148 & n7320 ;
  assign n7603 = x1146 & n7322 ;
  assign n7605 = n7604 ^ n7603 ;
  assign n7602 = n7307 ^ x273 ;
  assign n7606 = n7605 ^ n7602 ;
  assign n7601 = x1147 & ~n4095 ;
  assign n7607 = n7606 ^ n7601 ;
  assign n7608 = ~n7297 & n7607 ;
  assign n7609 = n7608 ^ n7602 ;
  assign n7615 = x1143 & n7322 ;
  assign n7614 = x1145 & n7320 ;
  assign n7616 = n7615 ^ n7614 ;
  assign n7611 = x659 ^ x274 ;
  assign n7612 = n7304 & ~n7611 ;
  assign n7613 = n7612 ^ x274 ;
  assign n7617 = n7616 ^ n7613 ;
  assign n7610 = x1144 & ~n4095 ;
  assign n7618 = n7617 ^ n7610 ;
  assign n7619 = ~n7297 & ~n7618 ;
  assign n7620 = n7619 ^ n7613 ;
  assign n7624 = x1149 & n7322 ;
  assign n7623 = x1151 & n7320 ;
  assign n7625 = n7624 ^ n7623 ;
  assign n7622 = n7310 ^ x275 ;
  assign n7626 = n7625 ^ n7622 ;
  assign n7621 = x1150 & ~n4095 ;
  assign n7627 = n7626 ^ n7621 ;
  assign n7628 = ~n7297 & n7627 ;
  assign n7629 = n7628 ^ n7622 ;
  assign n7633 = x1144 & n7322 ;
  assign n7632 = x1146 & n7320 ;
  assign n7634 = n7633 ^ n7632 ;
  assign n7631 = n7305 ^ x276 ;
  assign n7635 = n7634 ^ n7631 ;
  assign n7630 = x1145 & ~n4095 ;
  assign n7636 = n7635 ^ n7630 ;
  assign n7637 = ~n7297 & n7636 ;
  assign n7638 = n7637 ^ n7631 ;
  assign n7644 = x1142 & n7320 ;
  assign n7643 = x1140 & n7322 ;
  assign n7645 = n7644 ^ n7643 ;
  assign n7640 = x820 ^ x277 ;
  assign n7641 = n7304 & ~n7640 ;
  assign n7642 = n7641 ^ x277 ;
  assign n7646 = n7645 ^ n7642 ;
  assign n7639 = x1141 & ~n4095 ;
  assign n7647 = n7646 ^ n7639 ;
  assign n7648 = ~n7297 & ~n7647 ;
  assign n7649 = n7648 ^ n7642 ;
  assign n7657 = x1133 & ~n4095 ;
  assign n7655 = x1134 & n7320 ;
  assign n7653 = x1132 & n7322 ;
  assign n7650 = x976 ^ x278 ;
  assign n7651 = n7304 & n7650 ;
  assign n7652 = n7651 ^ x278 ;
  assign n7654 = n7653 ^ n7652 ;
  assign n7656 = n7655 ^ n7654 ;
  assign n7658 = n7657 ^ n7656 ;
  assign n7659 = ~n7297 & n7658 ;
  assign n7660 = n7659 ^ n7652 ;
  assign n7666 = x1135 & n7320 ;
  assign n7665 = x1133 & n7322 ;
  assign n7667 = n7666 ^ n7665 ;
  assign n7662 = x958 ^ x279 ;
  assign n7663 = n7304 & n7662 ;
  assign n7664 = n7663 ^ x279 ;
  assign n7668 = n7667 ^ n7664 ;
  assign n7661 = x1134 & ~n4095 ;
  assign n7669 = n7668 ^ n7661 ;
  assign n7670 = ~n7297 & n7669 ;
  assign n7671 = n7670 ^ n7664 ;
  assign n7677 = x1137 & n7320 ;
  assign n7676 = x1135 & n7322 ;
  assign n7678 = n7677 ^ n7676 ;
  assign n7673 = x914 ^ x280 ;
  assign n7674 = n7304 & ~n7673 ;
  assign n7675 = n7674 ^ x280 ;
  assign n7679 = n7678 ^ n7675 ;
  assign n7672 = x1136 & ~n4095 ;
  assign n7680 = n7679 ^ n7672 ;
  assign n7681 = ~n7297 & ~n7680 ;
  assign n7682 = n7681 ^ n7675 ;
  assign n7688 = x1139 & n7320 ;
  assign n7687 = x1137 & n7322 ;
  assign n7689 = n7688 ^ n7687 ;
  assign n7684 = x830 ^ x281 ;
  assign n7685 = n7304 & ~n7684 ;
  assign n7686 = n7685 ^ x281 ;
  assign n7690 = n7689 ^ n7686 ;
  assign n7683 = x1138 & ~n4095 ;
  assign n7691 = n7690 ^ n7683 ;
  assign n7692 = ~n7297 & ~n7691 ;
  assign n7693 = n7692 ^ n7686 ;
  assign n7699 = x1140 & n7320 ;
  assign n7698 = x1138 & n7322 ;
  assign n7700 = n7699 ^ n7698 ;
  assign n7695 = x836 ^ x282 ;
  assign n7696 = n7304 & ~n7695 ;
  assign n7697 = n7696 ^ x282 ;
  assign n7701 = n7700 ^ n7697 ;
  assign n7694 = x1139 & ~n4095 ;
  assign n7702 = n7701 ^ n7694 ;
  assign n7703 = ~n7297 & ~n7702 ;
  assign n7704 = n7703 ^ n7697 ;
  assign n7708 = x1147 & n7322 ;
  assign n7707 = x1149 & n7320 ;
  assign n7709 = n7708 ^ n7707 ;
  assign n7706 = n7308 ^ x283 ;
  assign n7710 = n7709 ^ n7706 ;
  assign n7705 = x1148 & ~n4095 ;
  assign n7711 = n7710 ^ n7705 ;
  assign n7712 = ~n7297 & n7711 ;
  assign n7713 = n7712 ^ n7706 ;
  assign n7720 = x1143 & n7014 ;
  assign n7721 = n4252 & n7720 ;
  assign n7722 = n7721 ^ n4252 ;
  assign n7714 = n4252 ^ x284 ;
  assign n7723 = n7722 ^ n7714 ;
  assign n7724 = ~n7492 & ~n7723 ;
  assign n7725 = n7724 ^ x284 ;
  assign n7726 = n4008 & n4215 ;
  assign n7727 = ~x288 & n3200 ;
  assign n7728 = ~n7726 & n7727 ;
  assign n7729 = x285 & n3197 ;
  assign n7730 = n7728 & n7729 ;
  assign n7733 = x286 & x288 ;
  assign n7736 = ~n3200 & n7726 ;
  assign n7745 = x288 & n7736 ;
  assign n7762 = n7733 & n7745 ;
  assign n7740 = x289 & n7762 ;
  assign n7741 = n7740 ^ x289 ;
  assign n7731 = x289 ^ x285 ;
  assign n7742 = n7741 ^ n7731 ;
  assign n7743 = ~x793 & n7742 ;
  assign n7744 = ~n7730 & n7743 ;
  assign n7746 = n7745 ^ x286 ;
  assign n7747 = n7746 ^ n7728 ;
  assign n7748 = ~x793 & n7747 ;
  assign n7750 = n3198 & n7748 ;
  assign n7751 = n7750 ^ n7748 ;
  assign n7752 = ~x287 & x457 ;
  assign n7753 = ~x332 & ~n7752 ;
  assign n7754 = n3201 ^ x288 ;
  assign n7755 = n7754 ^ n7726 ;
  assign n7756 = ~x793 & n7755 ;
  assign n7759 = ~x286 & n7728 ;
  assign n7760 = x289 & n7759 ;
  assign n7757 = n7730 ^ x289 ;
  assign n7761 = n7760 ^ n7757 ;
  assign n7763 = n7762 ^ n7761 ;
  assign n7764 = ~x793 & n7763 ;
  assign n7765 = x1048 ^ x290 ;
  assign n7766 = ~x476 & n7765 ;
  assign n7767 = n7766 ^ x290 ;
  assign n7768 = x1049 ^ x291 ;
  assign n7769 = ~x476 & n7768 ;
  assign n7770 = n7769 ^ x291 ;
  assign n7771 = x1084 ^ x292 ;
  assign n7772 = ~x476 & n7771 ;
  assign n7773 = n7772 ^ x292 ;
  assign n7774 = x1059 ^ x293 ;
  assign n7775 = ~x476 & n7774 ;
  assign n7776 = n7775 ^ x293 ;
  assign n7777 = x1072 ^ x294 ;
  assign n7778 = ~x476 & n7777 ;
  assign n7779 = n7778 ^ x294 ;
  assign n7780 = x1053 ^ x295 ;
  assign n7781 = ~x476 & n7780 ;
  assign n7782 = n7781 ^ x295 ;
  assign n7783 = x1037 ^ x296 ;
  assign n7784 = ~x476 & n7783 ;
  assign n7785 = n7784 ^ x296 ;
  assign n7786 = x1044 ^ x297 ;
  assign n7787 = ~x476 & n7786 ;
  assign n7788 = n7787 ^ x297 ;
  assign n7789 = x1044 ^ x298 ;
  assign n7790 = ~x478 & n7789 ;
  assign n7791 = n7790 ^ x298 ;
  assign n7797 = n1290 & n1323 ;
  assign n7792 = x39 & n3967 ;
  assign n7793 = ~x287 & n7792 ;
  assign n7794 = n7793 ^ n4258 ;
  assign n7796 = ~n4266 & ~n7794 ;
  assign n7799 = n7797 ^ n7796 ;
  assign n7800 = ~x24 & n1326 ;
  assign n7805 = ~x312 & n7800 ;
  assign n7806 = n7805 ^ x300 ;
  assign n7807 = ~x55 & ~n7806 ;
  assign n7808 = ~x300 & ~x312 ;
  assign n7813 = n7800 & n7808 ;
  assign n7814 = n7813 ^ x301 ;
  assign n7815 = ~x55 & ~n7814 ;
  assign n7820 = n2490 ^ n1916 ;
  assign n7821 = ~x237 & n7820 ;
  assign n7816 = n1931 ^ n1373 ;
  assign n7817 = n1537 & n7816 ;
  assign n7818 = n7817 ^ n1373 ;
  assign n7819 = x937 & n7818 ;
  assign n7822 = n7821 ^ n7819 ;
  assign n7827 = x1148 & n2588 ;
  assign n7823 = n1936 ^ n1350 ;
  assign n7824 = n1537 & n7823 ;
  assign n7825 = n7824 ^ n1350 ;
  assign n7826 = x273 & n7825 ;
  assign n7828 = n7827 ^ n7826 ;
  assign n7829 = ~n7822 & ~n7828 ;
  assign n7830 = x1049 ^ x303 ;
  assign n7831 = ~x478 & n7830 ;
  assign n7832 = n7831 ^ x303 ;
  assign n7833 = x1048 ^ x304 ;
  assign n7834 = ~x478 & n7833 ;
  assign n7835 = n7834 ^ x304 ;
  assign n7836 = x1084 ^ x305 ;
  assign n7837 = ~x478 & n7836 ;
  assign n7838 = n7837 ^ x305 ;
  assign n7839 = x1059 ^ x306 ;
  assign n7840 = ~x478 & n7839 ;
  assign n7841 = n7840 ^ x306 ;
  assign n7842 = x1053 ^ x307 ;
  assign n7843 = ~x478 & n7842 ;
  assign n7844 = n7843 ^ x307 ;
  assign n7845 = x1037 ^ x308 ;
  assign n7846 = ~x478 & n7845 ;
  assign n7847 = n7846 ^ x308 ;
  assign n7848 = x1072 ^ x309 ;
  assign n7849 = ~x478 & n7848 ;
  assign n7850 = n7849 ^ x309 ;
  assign n7852 = ~x233 & n7820 ;
  assign n7851 = x271 & n7825 ;
  assign n7853 = n7852 ^ n7851 ;
  assign n7855 = x934 & n7818 ;
  assign n7854 = x1147 & n2588 ;
  assign n7856 = n7855 ^ n7854 ;
  assign n7857 = ~n7853 & ~n7856 ;
  assign n7858 = x301 & n7808 ;
  assign n7863 = n7800 & n7858 ;
  assign n7864 = n7863 ^ x311 ;
  assign n7865 = ~x55 & ~n7864 ;
  assign n7866 = n7800 ^ x312 ;
  assign n7867 = ~x55 & n7866 ;
  assign n7868 = n4899 ^ n2608 ;
  assign n7869 = n4885 ^ x314 ;
  assign n7872 = ~n4899 & n7869 ;
  assign n7873 = n7872 ^ x314 ;
  assign n7874 = n7868 & ~n7873 ;
  assign n7875 = n7874 ^ n2608 ;
  assign n7876 = n7875 ^ x313 ;
  assign n7877 = ~x954 & ~n7876 ;
  assign n7878 = n7877 ^ x313 ;
  assign n7879 = n5154 & n5444 ;
  assign n7880 = ~x340 & n7726 ;
  assign n7881 = x1080 ^ x315 ;
  assign n7882 = n7880 & n7881 ;
  assign n7883 = n7882 ^ x315 ;
  assign n7884 = x1047 ^ x316 ;
  assign n7885 = n7880 & n7884 ;
  assign n7886 = n7885 ^ x316 ;
  assign n7887 = ~x330 & n7726 ;
  assign n7888 = x1078 ^ x317 ;
  assign n7889 = n7887 & n7888 ;
  assign n7890 = n7889 ^ x317 ;
  assign n7891 = ~x341 & n7726 ;
  assign n7892 = x1074 ^ x318 ;
  assign n7893 = n7891 & n7892 ;
  assign n7894 = n7893 ^ x318 ;
  assign n7895 = x1072 ^ x319 ;
  assign n7896 = n7891 & n7895 ;
  assign n7897 = n7896 ^ x319 ;
  assign n7898 = x1048 ^ x320 ;
  assign n7899 = n7880 & n7898 ;
  assign n7900 = n7899 ^ x320 ;
  assign n7901 = x1058 ^ x321 ;
  assign n7902 = n7880 & n7901 ;
  assign n7903 = n7902 ^ x321 ;
  assign n7904 = x1051 ^ x322 ;
  assign n7905 = n7880 & n7904 ;
  assign n7906 = n7905 ^ x322 ;
  assign n7907 = x1065 ^ x323 ;
  assign n7908 = n7880 & n7907 ;
  assign n7909 = n7908 ^ x323 ;
  assign n7910 = x1086 ^ x324 ;
  assign n7911 = n7891 & n7910 ;
  assign n7912 = n7911 ^ x324 ;
  assign n7913 = x1063 ^ x325 ;
  assign n7914 = n7891 & n7913 ;
  assign n7915 = n7914 ^ x325 ;
  assign n7916 = x1057 ^ x326 ;
  assign n7917 = n7891 & n7916 ;
  assign n7918 = n7917 ^ x326 ;
  assign n7919 = x1040 ^ x327 ;
  assign n7920 = n7880 & n7919 ;
  assign n7921 = n7920 ^ x327 ;
  assign n7922 = x1058 ^ x328 ;
  assign n7923 = n7891 & n7922 ;
  assign n7924 = n7923 ^ x328 ;
  assign n7925 = x1043 ^ x329 ;
  assign n7926 = n7891 & n7925 ;
  assign n7927 = n7926 ^ x329 ;
  assign n7928 = x1091 & n3009 ;
  assign n7929 = n7928 ^ x1092 ;
  assign n7930 = n7887 ^ n7880 ;
  assign n7931 = n7930 ^ x330 ;
  assign n7932 = n7929 & ~n7931 ;
  assign n7934 = ~x331 & n7726 ;
  assign n7933 = n7891 ^ x331 ;
  assign n7935 = n7934 ^ n7933 ;
  assign n7936 = n7929 & ~n7935 ;
  assign n7939 = n1919 & n3934 ;
  assign n7937 = ~n1309 & ~n3964 ;
  assign n7938 = ~n4129 & n7937 ;
  assign n7941 = n7939 ^ n7938 ;
  assign n7942 = x1040 ^ x333 ;
  assign n7943 = n7891 & n7942 ;
  assign n7944 = n7943 ^ x333 ;
  assign n7945 = x1065 ^ x334 ;
  assign n7946 = n7891 & n7945 ;
  assign n7947 = n7946 ^ x334 ;
  assign n7948 = x1069 ^ x335 ;
  assign n7949 = n7891 & n7948 ;
  assign n7950 = n7949 ^ x335 ;
  assign n7951 = x1070 ^ x336 ;
  assign n7952 = n7887 & n7951 ;
  assign n7953 = n7952 ^ x336 ;
  assign n7954 = x1044 ^ x337 ;
  assign n7955 = n7887 & n7954 ;
  assign n7956 = n7955 ^ x337 ;
  assign n7957 = x1072 ^ x338 ;
  assign n7958 = n7887 & n7957 ;
  assign n7959 = n7958 ^ x338 ;
  assign n7960 = x1086 ^ x339 ;
  assign n7961 = n7887 & n7960 ;
  assign n7962 = n7961 ^ x339 ;
  assign n7963 = n7880 ^ x340 ;
  assign n7964 = n7963 ^ n7934 ;
  assign n7965 = n7929 & n7964 ;
  assign n7966 = n7891 ^ n7887 ;
  assign n7967 = n7966 ^ x341 ;
  assign n7968 = n7929 & ~n7967 ;
  assign n7969 = x1049 ^ x342 ;
  assign n7970 = n7880 & n7969 ;
  assign n7971 = n7970 ^ x342 ;
  assign n7972 = x1062 ^ x343 ;
  assign n7973 = n7880 & n7972 ;
  assign n7974 = n7973 ^ x343 ;
  assign n7975 = x1069 ^ x344 ;
  assign n7976 = n7880 & n7975 ;
  assign n7977 = n7976 ^ x344 ;
  assign n7978 = x1039 ^ x345 ;
  assign n7979 = n7880 & n7978 ;
  assign n7980 = n7979 ^ x345 ;
  assign n7981 = x1067 ^ x346 ;
  assign n7982 = n7880 & n7981 ;
  assign n7983 = n7982 ^ x346 ;
  assign n7984 = x1055 ^ x347 ;
  assign n7985 = n7880 & n7984 ;
  assign n7986 = n7985 ^ x347 ;
  assign n7987 = x1087 ^ x348 ;
  assign n7988 = n7880 & n7987 ;
  assign n7989 = n7988 ^ x348 ;
  assign n7990 = x1043 ^ x349 ;
  assign n7991 = n7880 & n7990 ;
  assign n7992 = n7991 ^ x349 ;
  assign n7993 = x1035 ^ x350 ;
  assign n7994 = n7880 & n7993 ;
  assign n7995 = n7994 ^ x350 ;
  assign n7996 = x1079 ^ x351 ;
  assign n7997 = n7880 & n7996 ;
  assign n7998 = n7997 ^ x351 ;
  assign n7999 = x1078 ^ x352 ;
  assign n8000 = n7880 & n7999 ;
  assign n8001 = n8000 ^ x352 ;
  assign n8002 = x1063 ^ x353 ;
  assign n8003 = n7880 & n8002 ;
  assign n8004 = n8003 ^ x353 ;
  assign n8005 = x1045 ^ x354 ;
  assign n8006 = n7880 & n8005 ;
  assign n8007 = n8006 ^ x354 ;
  assign n8008 = x1084 ^ x355 ;
  assign n8009 = n7880 & n8008 ;
  assign n8010 = n8009 ^ x355 ;
  assign n8011 = x1081 ^ x356 ;
  assign n8012 = n7880 & n8011 ;
  assign n8013 = n8012 ^ x356 ;
  assign n8014 = x1076 ^ x357 ;
  assign n8015 = n7880 & n8014 ;
  assign n8016 = n8015 ^ x357 ;
  assign n8017 = x1071 ^ x358 ;
  assign n8018 = n7880 & n8017 ;
  assign n8019 = n8018 ^ x358 ;
  assign n8020 = x1068 ^ x359 ;
  assign n8021 = n7880 & n8020 ;
  assign n8022 = n8021 ^ x359 ;
  assign n8023 = x1042 ^ x360 ;
  assign n8024 = n7880 & n8023 ;
  assign n8025 = n8024 ^ x360 ;
  assign n8026 = x1059 ^ x361 ;
  assign n8027 = n7880 & n8026 ;
  assign n8028 = n8027 ^ x361 ;
  assign n8029 = x1070 ^ x362 ;
  assign n8030 = n7880 & n8029 ;
  assign n8031 = n8030 ^ x362 ;
  assign n8032 = x1049 ^ x363 ;
  assign n8033 = n7887 & n8032 ;
  assign n8034 = n8033 ^ x363 ;
  assign n8035 = x1062 ^ x364 ;
  assign n8036 = n7887 & n8035 ;
  assign n8037 = n8036 ^ x364 ;
  assign n8038 = x1065 ^ x365 ;
  assign n8039 = n7887 & n8038 ;
  assign n8040 = n8039 ^ x365 ;
  assign n8041 = x1069 ^ x366 ;
  assign n8042 = n7887 & n8041 ;
  assign n8043 = n8042 ^ x366 ;
  assign n8044 = x1039 ^ x367 ;
  assign n8045 = n7887 & n8044 ;
  assign n8046 = n8045 ^ x367 ;
  assign n8047 = x1067 ^ x368 ;
  assign n8048 = n7887 & n8047 ;
  assign n8049 = n8048 ^ x368 ;
  assign n8050 = x1080 ^ x369 ;
  assign n8051 = n7887 & n8050 ;
  assign n8052 = n8051 ^ x369 ;
  assign n8053 = x1055 ^ x370 ;
  assign n8054 = n7887 & n8053 ;
  assign n8055 = n8054 ^ x370 ;
  assign n8056 = x1051 ^ x371 ;
  assign n8057 = n7887 & n8056 ;
  assign n8058 = n8057 ^ x371 ;
  assign n8059 = x1048 ^ x372 ;
  assign n8060 = n7887 & n8059 ;
  assign n8061 = n8060 ^ x372 ;
  assign n8062 = x1087 ^ x373 ;
  assign n8063 = n7887 & n8062 ;
  assign n8064 = n8063 ^ x373 ;
  assign n8065 = x1035 ^ x374 ;
  assign n8066 = n7887 & n8065 ;
  assign n8067 = n8066 ^ x374 ;
  assign n8068 = x1047 ^ x375 ;
  assign n8069 = n7887 & n8068 ;
  assign n8070 = n8069 ^ x375 ;
  assign n8071 = x1079 ^ x376 ;
  assign n8072 = n7887 & n8071 ;
  assign n8073 = n8072 ^ x376 ;
  assign n8074 = x1074 ^ x377 ;
  assign n8075 = n7887 & n8074 ;
  assign n8076 = n8075 ^ x377 ;
  assign n8077 = x1063 ^ x378 ;
  assign n8078 = n7887 & n8077 ;
  assign n8079 = n8078 ^ x378 ;
  assign n8080 = x1045 ^ x379 ;
  assign n8081 = n7887 & n8080 ;
  assign n8082 = n8081 ^ x379 ;
  assign n8083 = x1084 ^ x380 ;
  assign n8084 = n7887 & n8083 ;
  assign n8085 = n8084 ^ x380 ;
  assign n8086 = x1081 ^ x381 ;
  assign n8087 = n7887 & n8086 ;
  assign n8088 = n8087 ^ x381 ;
  assign n8089 = x1076 ^ x382 ;
  assign n8090 = n7887 & n8089 ;
  assign n8091 = n8090 ^ x382 ;
  assign n8092 = x1071 ^ x383 ;
  assign n8093 = n7887 & n8092 ;
  assign n8094 = n8093 ^ x383 ;
  assign n8095 = x1068 ^ x384 ;
  assign n8096 = n7887 & n8095 ;
  assign n8097 = n8096 ^ x384 ;
  assign n8098 = x1042 ^ x385 ;
  assign n8099 = n7887 & n8098 ;
  assign n8100 = n8099 ^ x385 ;
  assign n8101 = x1059 ^ x386 ;
  assign n8102 = n7887 & n8101 ;
  assign n8103 = n8102 ^ x386 ;
  assign n8104 = x1053 ^ x387 ;
  assign n8105 = n7887 & n8104 ;
  assign n8106 = n8105 ^ x387 ;
  assign n8107 = x1037 ^ x388 ;
  assign n8108 = n7887 & n8107 ;
  assign n8109 = n8108 ^ x388 ;
  assign n8110 = x1036 ^ x389 ;
  assign n8111 = n7887 & n8110 ;
  assign n8112 = n8111 ^ x389 ;
  assign n8113 = x1049 ^ x390 ;
  assign n8114 = n7891 & n8113 ;
  assign n8115 = n8114 ^ x390 ;
  assign n8116 = x1062 ^ x391 ;
  assign n8117 = n7891 & n8116 ;
  assign n8118 = n8117 ^ x391 ;
  assign n8119 = x1039 ^ x392 ;
  assign n8120 = n7891 & n8119 ;
  assign n8121 = n8120 ^ x392 ;
  assign n8122 = x1067 ^ x393 ;
  assign n8123 = n7891 & n8122 ;
  assign n8124 = n8123 ^ x393 ;
  assign n8125 = x1080 ^ x394 ;
  assign n8126 = n7891 & n8125 ;
  assign n8127 = n8126 ^ x394 ;
  assign n8128 = x1055 ^ x395 ;
  assign n8129 = n7891 & n8128 ;
  assign n8130 = n8129 ^ x395 ;
  assign n8131 = x1051 ^ x396 ;
  assign n8132 = n7891 & n8131 ;
  assign n8133 = n8132 ^ x396 ;
  assign n8134 = x1048 ^ x397 ;
  assign n8135 = n7891 & n8134 ;
  assign n8136 = n8135 ^ x397 ;
  assign n8137 = x1087 ^ x398 ;
  assign n8138 = n7891 & n8137 ;
  assign n8139 = n8138 ^ x398 ;
  assign n8140 = x1047 ^ x399 ;
  assign n8141 = n7891 & n8140 ;
  assign n8142 = n8141 ^ x399 ;
  assign n8143 = x1035 ^ x400 ;
  assign n8144 = n7891 & n8143 ;
  assign n8145 = n8144 ^ x400 ;
  assign n8146 = x1079 ^ x401 ;
  assign n8147 = n7891 & n8146 ;
  assign n8148 = n8147 ^ x401 ;
  assign n8149 = x1078 ^ x402 ;
  assign n8150 = n7891 & n8149 ;
  assign n8151 = n8150 ^ x402 ;
  assign n8152 = x1045 ^ x403 ;
  assign n8153 = n7891 & n8152 ;
  assign n8154 = n8153 ^ x403 ;
  assign n8155 = x1084 ^ x404 ;
  assign n8156 = n7891 & n8155 ;
  assign n8157 = n8156 ^ x404 ;
  assign n8158 = x1081 ^ x405 ;
  assign n8159 = n7891 & n8158 ;
  assign n8160 = n8159 ^ x405 ;
  assign n8161 = x1076 ^ x406 ;
  assign n8162 = n7891 & n8161 ;
  assign n8163 = n8162 ^ x406 ;
  assign n8164 = x1071 ^ x407 ;
  assign n8165 = n7891 & n8164 ;
  assign n8166 = n8165 ^ x407 ;
  assign n8167 = x1068 ^ x408 ;
  assign n8168 = n7891 & n8167 ;
  assign n8169 = n8168 ^ x408 ;
  assign n8170 = x1042 ^ x409 ;
  assign n8171 = n7891 & n8170 ;
  assign n8172 = n8171 ^ x409 ;
  assign n8173 = x1059 ^ x410 ;
  assign n8174 = n7891 & n8173 ;
  assign n8175 = n8174 ^ x410 ;
  assign n8176 = x1053 ^ x411 ;
  assign n8177 = n7891 & n8176 ;
  assign n8178 = n8177 ^ x411 ;
  assign n8179 = x1037 ^ x412 ;
  assign n8180 = n7891 & n8179 ;
  assign n8181 = n8180 ^ x412 ;
  assign n8182 = x1036 ^ x413 ;
  assign n8183 = n7891 & n8182 ;
  assign n8184 = n8183 ^ x413 ;
  assign n8185 = x1049 ^ x414 ;
  assign n8186 = n7934 & n8185 ;
  assign n8187 = n8186 ^ x414 ;
  assign n8188 = x1062 ^ x415 ;
  assign n8189 = n7934 & n8188 ;
  assign n8190 = n8189 ^ x415 ;
  assign n8191 = x1069 ^ x416 ;
  assign n8192 = n7934 & n8191 ;
  assign n8193 = n8192 ^ x416 ;
  assign n8194 = x1039 ^ x417 ;
  assign n8195 = n7934 & n8194 ;
  assign n8196 = n8195 ^ x417 ;
  assign n8197 = x1067 ^ x418 ;
  assign n8198 = n7934 & n8197 ;
  assign n8199 = n8198 ^ x418 ;
  assign n8200 = x1080 ^ x419 ;
  assign n8201 = n7934 & n8200 ;
  assign n8202 = n8201 ^ x419 ;
  assign n8203 = x1055 ^ x420 ;
  assign n8204 = n7934 & n8203 ;
  assign n8205 = n8204 ^ x420 ;
  assign n8206 = x1051 ^ x421 ;
  assign n8207 = n7934 & n8206 ;
  assign n8208 = n8207 ^ x421 ;
  assign n8209 = x1048 ^ x422 ;
  assign n8210 = n7934 & n8209 ;
  assign n8211 = n8210 ^ x422 ;
  assign n8212 = x1087 ^ x423 ;
  assign n8213 = n7934 & n8212 ;
  assign n8214 = n8213 ^ x423 ;
  assign n8215 = x1047 ^ x424 ;
  assign n8216 = n7934 & n8215 ;
  assign n8217 = n8216 ^ x424 ;
  assign n8218 = x1035 ^ x425 ;
  assign n8219 = n7934 & n8218 ;
  assign n8220 = n8219 ^ x425 ;
  assign n8221 = x1079 ^ x426 ;
  assign n8222 = n7934 & n8221 ;
  assign n8223 = n8222 ^ x426 ;
  assign n8224 = x1078 ^ x427 ;
  assign n8225 = n7934 & n8224 ;
  assign n8226 = n8225 ^ x427 ;
  assign n8227 = x1045 ^ x428 ;
  assign n8228 = n7934 & n8227 ;
  assign n8229 = n8228 ^ x428 ;
  assign n8230 = x1084 ^ x429 ;
  assign n8231 = n7934 & n8230 ;
  assign n8232 = n8231 ^ x429 ;
  assign n8233 = x1076 ^ x430 ;
  assign n8234 = n7934 & n8233 ;
  assign n8235 = n8234 ^ x430 ;
  assign n8236 = x1071 ^ x431 ;
  assign n8237 = n7934 & n8236 ;
  assign n8238 = n8237 ^ x431 ;
  assign n8239 = x1068 ^ x432 ;
  assign n8240 = n7934 & n8239 ;
  assign n8241 = n8240 ^ x432 ;
  assign n8242 = x1042 ^ x433 ;
  assign n8243 = n7934 & n8242 ;
  assign n8244 = n8243 ^ x433 ;
  assign n8245 = x1059 ^ x434 ;
  assign n8246 = n7934 & n8245 ;
  assign n8247 = n8246 ^ x434 ;
  assign n8248 = x1053 ^ x435 ;
  assign n8249 = n7934 & n8248 ;
  assign n8250 = n8249 ^ x435 ;
  assign n8251 = x1037 ^ x436 ;
  assign n8252 = n7934 & n8251 ;
  assign n8253 = n8252 ^ x436 ;
  assign n8254 = x1070 ^ x437 ;
  assign n8255 = n7934 & n8254 ;
  assign n8256 = n8255 ^ x437 ;
  assign n8257 = x1036 ^ x438 ;
  assign n8258 = n7934 & n8257 ;
  assign n8259 = n8258 ^ x438 ;
  assign n8260 = x1057 ^ x439 ;
  assign n8261 = n7887 & n8260 ;
  assign n8262 = n8261 ^ x439 ;
  assign n8263 = x1043 ^ x440 ;
  assign n8264 = n7887 & n8263 ;
  assign n8265 = n8264 ^ x440 ;
  assign n8266 = x1044 ^ x441 ;
  assign n8267 = n7880 & n8266 ;
  assign n8268 = n8267 ^ x441 ;
  assign n8269 = x1058 ^ x442 ;
  assign n8270 = n7887 & n8269 ;
  assign n8271 = n8270 ^ x442 ;
  assign n8272 = x1044 ^ x443 ;
  assign n8273 = n7934 & n8272 ;
  assign n8274 = n8273 ^ x443 ;
  assign n8275 = x1072 ^ x444 ;
  assign n8276 = n7934 & n8275 ;
  assign n8277 = n8276 ^ x444 ;
  assign n8278 = x1081 ^ x445 ;
  assign n8279 = n7934 & n8278 ;
  assign n8280 = n8279 ^ x445 ;
  assign n8281 = x1086 ^ x446 ;
  assign n8282 = n7934 & n8281 ;
  assign n8283 = n8282 ^ x446 ;
  assign n8284 = x1040 ^ x447 ;
  assign n8285 = n7887 & n8284 ;
  assign n8286 = n8285 ^ x447 ;
  assign n8287 = x1074 ^ x448 ;
  assign n8288 = n7934 & n8287 ;
  assign n8289 = n8288 ^ x448 ;
  assign n8290 = x1057 ^ x449 ;
  assign n8291 = n7934 & n8290 ;
  assign n8292 = n8291 ^ x449 ;
  assign n8293 = x1036 ^ x450 ;
  assign n8294 = n7880 & n8293 ;
  assign n8295 = n8294 ^ x450 ;
  assign n8296 = x1063 ^ x451 ;
  assign n8297 = n7934 & n8296 ;
  assign n8298 = n8297 ^ x451 ;
  assign n8299 = x1053 ^ x452 ;
  assign n8300 = n7880 & n8299 ;
  assign n8301 = n8300 ^ x452 ;
  assign n8302 = x1040 ^ x453 ;
  assign n8303 = n7934 & n8302 ;
  assign n8304 = n8303 ^ x453 ;
  assign n8305 = x1043 ^ x454 ;
  assign n8306 = n7934 & n8305 ;
  assign n8307 = n8306 ^ x454 ;
  assign n8308 = x1037 ^ x455 ;
  assign n8309 = n7880 & n8308 ;
  assign n8310 = n8309 ^ x455 ;
  assign n8311 = x1044 ^ x456 ;
  assign n8312 = n7891 & n8311 ;
  assign n8313 = n8312 ^ x456 ;
  assign n8314 = x594 & x600 ;
  assign n8315 = x597 & x601 ;
  assign n8316 = n8314 & n8315 ;
  assign n8317 = n8316 ^ x804 ;
  assign n8318 = n8317 ^ x595 ;
  assign n8321 = x804 ^ x596 ;
  assign n8322 = n8321 ^ x810 ;
  assign n8323 = x815 ^ x804 ;
  assign n8324 = n8323 ^ n8322 ;
  assign n8325 = x815 ^ x810 ;
  assign n8326 = n8325 ^ n8322 ;
  assign n8327 = x810 ^ x599 ;
  assign n8328 = n8327 ^ x804 ;
  assign n8329 = n8326 & n8328 ;
  assign n8330 = n8324 & n8329 ;
  assign n8331 = n8330 ^ x810 ;
  assign n8332 = n8331 ^ x804 ;
  assign n8333 = n8322 & n8332 ;
  assign n8334 = x804 & n8333 ;
  assign n8319 = x810 ^ x804 ;
  assign n8335 = n8334 ^ n8319 ;
  assign n8336 = n8318 & n8335 ;
  assign n8337 = n8336 ^ x804 ;
  assign n8338 = n8316 & ~n8337 ;
  assign n8339 = x600 & x804 ;
  assign n8340 = ~x810 & n8339 ;
  assign n8341 = n8340 ^ x804 ;
  assign n8342 = ~x601 & ~x815 ;
  assign n8350 = ~x804 & n8342 ;
  assign n8351 = ~x810 & n8350 ;
  assign n8352 = n8351 ^ x810 ;
  assign n8343 = n8342 ^ x815 ;
  assign n8344 = n8343 ^ x810 ;
  assign n8353 = n8352 ^ n8344 ;
  assign n8354 = ~n8341 & ~n8353 ;
  assign n8355 = ~n8338 & ~n8354 ;
  assign n8356 = x605 & ~n8355 ;
  assign n8357 = ~x815 & x990 ;
  assign n8358 = n8314 & n8341 ;
  assign n8359 = n8357 & n8358 ;
  assign n8360 = ~n8356 & ~n8359 ;
  assign n8361 = x821 & ~n8360 ;
  assign n8362 = x1072 ^ x458 ;
  assign n8363 = n7880 & n8362 ;
  assign n8364 = n8363 ^ x458 ;
  assign n8365 = x1058 ^ x459 ;
  assign n8366 = n7934 & n8365 ;
  assign n8367 = n8366 ^ x459 ;
  assign n8368 = x1086 ^ x460 ;
  assign n8369 = n7880 & n8368 ;
  assign n8370 = n8369 ^ x460 ;
  assign n8371 = x1057 ^ x461 ;
  assign n8372 = n7880 & n8371 ;
  assign n8373 = n8372 ^ x461 ;
  assign n8374 = x1074 ^ x462 ;
  assign n8375 = n7880 & n8374 ;
  assign n8376 = n8375 ^ x462 ;
  assign n8377 = x1070 ^ x463 ;
  assign n8378 = n7891 & n8377 ;
  assign n8379 = n8378 ^ x463 ;
  assign n8380 = x1065 ^ x464 ;
  assign n8381 = n7934 & n8380 ;
  assign n8382 = n8381 ^ x464 ;
  assign n8385 = x1157 & n2588 ;
  assign n8384 = ~x243 & n7825 ;
  assign n8386 = n8385 ^ n8384 ;
  assign n8383 = x926 & n7818 ;
  assign n8387 = n8386 ^ n8383 ;
  assign n8390 = x1151 & n2588 ;
  assign n8389 = x275 & n7825 ;
  assign n8391 = n8390 ^ n8389 ;
  assign n8388 = x943 & n7818 ;
  assign n8392 = n8391 ^ n8388 ;
  assign n8394 = x40 & x1001 ;
  assign n8395 = n2650 & n2698 ;
  assign n8396 = n8394 & n8395 ;
  assign n8393 = n4325 & n6811 ;
  assign n8398 = n8396 ^ n8393 ;
  assign n8399 = x468 & ~n3943 ;
  assign n8400 = ~n4299 & n8399 ;
  assign n8401 = n8400 ^ n4299 ;
  assign n8404 = x1156 & n2588 ;
  assign n8403 = ~x263 & n7825 ;
  assign n8405 = n8404 ^ n8403 ;
  assign n8402 = x942 & n7818 ;
  assign n8406 = n8405 ^ n8402 ;
  assign n8409 = x1155 & n2588 ;
  assign n8408 = x267 & n7825 ;
  assign n8410 = n8409 ^ n8408 ;
  assign n8407 = x925 & n7818 ;
  assign n8411 = n8410 ^ n8407 ;
  assign n8414 = x1153 & n2588 ;
  assign n8413 = x253 & n7825 ;
  assign n8415 = n8414 ^ n8413 ;
  assign n8412 = x941 & n7818 ;
  assign n8416 = n8415 ^ n8412 ;
  assign n8419 = x1154 & n2588 ;
  assign n8418 = x254 & n7825 ;
  assign n8420 = n8419 ^ n8418 ;
  assign n8417 = x923 & n7818 ;
  assign n8421 = n8420 ^ n8417 ;
  assign n8424 = x1152 & n2588 ;
  assign n8423 = x268 & n7825 ;
  assign n8425 = n8424 ^ n8423 ;
  assign n8422 = x922 & n7818 ;
  assign n8426 = n8425 ^ n8422 ;
  assign n8429 = x1150 & n2588 ;
  assign n8428 = x272 & n7825 ;
  assign n8430 = n8429 ^ n8428 ;
  assign n8427 = x931 & n7818 ;
  assign n8431 = n8430 ^ n8427 ;
  assign n8434 = x1149 & n2588 ;
  assign n8433 = x283 & n7825 ;
  assign n8435 = n8434 ^ n8433 ;
  assign n8432 = x936 & n7818 ;
  assign n8436 = n8435 ^ n8432 ;
  assign n8437 = x71 & ~n4095 ;
  assign n8439 = n8437 ^ n4652 ;
  assign n8440 = x71 & n7322 ;
  assign n8441 = x481 ^ x248 ;
  assign n8442 = ~n6508 & n8441 ;
  assign n8443 = n8442 ^ x248 ;
  assign n8444 = x482 ^ x249 ;
  assign n8445 = ~n6524 & n8444 ;
  assign n8446 = n8445 ^ x249 ;
  assign n8447 = x483 ^ x242 ;
  assign n8448 = ~n6556 & n8447 ;
  assign n8449 = n8448 ^ x242 ;
  assign n8450 = x484 ^ x249 ;
  assign n8451 = ~n6556 & n8450 ;
  assign n8452 = n8451 ^ x249 ;
  assign n8453 = x485 ^ x234 ;
  assign n8454 = ~n6555 & n8453 ;
  assign n8455 = n8454 ^ x234 ;
  assign n8456 = x486 ^ x244 ;
  assign n8457 = ~n6555 & n8456 ;
  assign n8458 = n8457 ^ x244 ;
  assign n8459 = x487 ^ x246 ;
  assign n8460 = ~n6508 & n8459 ;
  assign n8461 = n8460 ^ x246 ;
  assign n8462 = x488 ^ x239 ;
  assign n8463 = ~n6508 & ~n8462 ;
  assign n8464 = n8463 ^ x239 ;
  assign n8465 = x489 ^ x242 ;
  assign n8466 = ~n6555 & n8465 ;
  assign n8467 = n8466 ^ x242 ;
  assign n8468 = x490 ^ x241 ;
  assign n8469 = ~n6556 & n8468 ;
  assign n8470 = n8469 ^ x241 ;
  assign n8471 = x491 ^ x238 ;
  assign n8472 = ~n6556 & n8471 ;
  assign n8473 = n8472 ^ x238 ;
  assign n8474 = x492 ^ x240 ;
  assign n8475 = ~n6556 & n8474 ;
  assign n8476 = n8475 ^ x240 ;
  assign n8477 = x493 ^ x244 ;
  assign n8478 = ~n6556 & n8477 ;
  assign n8479 = n8478 ^ x244 ;
  assign n8480 = x494 ^ x239 ;
  assign n8481 = ~n6556 & ~n8480 ;
  assign n8482 = n8481 ^ x239 ;
  assign n8483 = x495 ^ x235 ;
  assign n8484 = ~n6556 & n8483 ;
  assign n8485 = n8484 ^ x235 ;
  assign n8486 = x496 ^ x249 ;
  assign n8487 = ~n6541 & n8486 ;
  assign n8488 = n8487 ^ x249 ;
  assign n8489 = x497 ^ x239 ;
  assign n8490 = ~n6541 & ~n8489 ;
  assign n8491 = n8490 ^ x239 ;
  assign n8492 = x498 ^ x238 ;
  assign n8493 = ~n6524 & n8492 ;
  assign n8494 = n8493 ^ x238 ;
  assign n8495 = x499 ^ x246 ;
  assign n8496 = ~n6541 & n8495 ;
  assign n8497 = n8496 ^ x246 ;
  assign n8498 = x500 ^ x241 ;
  assign n8499 = ~n6541 & n8498 ;
  assign n8500 = n8499 ^ x241 ;
  assign n8501 = x501 ^ x248 ;
  assign n8502 = ~n6541 & n8501 ;
  assign n8503 = n8502 ^ x248 ;
  assign n8504 = x502 ^ x247 ;
  assign n8505 = ~n6541 & n8504 ;
  assign n8506 = n8505 ^ x247 ;
  assign n8507 = x503 ^ x245 ;
  assign n8508 = ~n6541 & n8507 ;
  assign n8509 = n8508 ^ x245 ;
  assign n8510 = x504 ^ x242 ;
  assign n8511 = ~n6542 & n8510 ;
  assign n8512 = n8511 ^ x242 ;
  assign n8513 = x505 ^ x234 ;
  assign n8514 = ~n6541 & n8513 ;
  assign n8515 = n8514 ^ x234 ;
  assign n8516 = x506 ^ x241 ;
  assign n8517 = ~n6542 & n8516 ;
  assign n8518 = n8517 ^ x241 ;
  assign n8519 = x507 ^ x238 ;
  assign n8520 = ~n6542 & n8519 ;
  assign n8521 = n8520 ^ x238 ;
  assign n8522 = x508 ^ x247 ;
  assign n8523 = ~n6542 & n8522 ;
  assign n8524 = n8523 ^ x247 ;
  assign n8525 = x509 ^ x245 ;
  assign n8526 = ~n6542 & n8525 ;
  assign n8527 = n8526 ^ x245 ;
  assign n8528 = x510 ^ x242 ;
  assign n8529 = ~n6508 & n8528 ;
  assign n8530 = n8529 ^ x242 ;
  assign n8531 = x511 ^ x234 ;
  assign n8532 = ~n6508 & n8531 ;
  assign n8533 = n8532 ^ x234 ;
  assign n8534 = x512 ^ x235 ;
  assign n8535 = ~n6508 & n8534 ;
  assign n8536 = n8535 ^ x235 ;
  assign n8537 = x513 ^ x244 ;
  assign n8538 = ~n6508 & n8537 ;
  assign n8539 = n8538 ^ x244 ;
  assign n8540 = x514 ^ x245 ;
  assign n8541 = ~n6508 & n8540 ;
  assign n8542 = n8541 ^ x245 ;
  assign n8543 = x515 ^ x240 ;
  assign n8544 = ~n6508 & n8543 ;
  assign n8545 = n8544 ^ x240 ;
  assign n8546 = x516 ^ x247 ;
  assign n8547 = ~n6508 & n8546 ;
  assign n8548 = n8547 ^ x247 ;
  assign n8549 = x517 ^ x238 ;
  assign n8550 = ~n6508 & n8549 ;
  assign n8551 = n8550 ^ x238 ;
  assign n8552 = x518 ^ x234 ;
  assign n8553 = ~n6517 & n8552 ;
  assign n8554 = n8553 ^ x234 ;
  assign n8555 = x519 ^ x239 ;
  assign n8556 = ~n6517 & ~n8555 ;
  assign n8557 = n8556 ^ x239 ;
  assign n8558 = x520 ^ x246 ;
  assign n8559 = ~n6517 & n8558 ;
  assign n8560 = n8559 ^ x246 ;
  assign n8561 = x521 ^ x248 ;
  assign n8562 = ~n6517 & n8561 ;
  assign n8563 = n8562 ^ x248 ;
  assign n8564 = x522 ^ x238 ;
  assign n8565 = ~n6517 & n8564 ;
  assign n8566 = n8565 ^ x238 ;
  assign n8567 = x523 ^ x234 ;
  assign n8568 = ~n6690 & n8567 ;
  assign n8569 = n8568 ^ x234 ;
  assign n8570 = x524 ^ x239 ;
  assign n8571 = ~n6690 & ~n8570 ;
  assign n8572 = n8571 ^ x239 ;
  assign n8573 = x525 ^ x245 ;
  assign n8574 = ~n6690 & n8573 ;
  assign n8575 = n8574 ^ x245 ;
  assign n8576 = x526 ^ x246 ;
  assign n8577 = ~n6690 & n8576 ;
  assign n8578 = n8577 ^ x246 ;
  assign n8579 = x527 ^ x247 ;
  assign n8580 = ~n6690 & n8579 ;
  assign n8581 = n8580 ^ x247 ;
  assign n8582 = x528 ^ x249 ;
  assign n8583 = ~n6690 & n8582 ;
  assign n8584 = n8583 ^ x249 ;
  assign n8585 = x529 ^ x238 ;
  assign n8586 = ~n6690 & n8585 ;
  assign n8587 = n8586 ^ x238 ;
  assign n8588 = x530 ^ x240 ;
  assign n8589 = ~n6690 & n8588 ;
  assign n8590 = n8589 ^ x240 ;
  assign n8591 = x531 ^ x235 ;
  assign n8592 = ~n6524 & n8591 ;
  assign n8593 = n8592 ^ x235 ;
  assign n8594 = x532 ^ x247 ;
  assign n8595 = ~n6524 & n8594 ;
  assign n8596 = n8595 ^ x247 ;
  assign n8597 = x533 ^ x235 ;
  assign n8598 = ~n6542 & n8597 ;
  assign n8599 = n8598 ^ x235 ;
  assign n8600 = x534 ^ x239 ;
  assign n8601 = ~n6542 & ~n8600 ;
  assign n8602 = n8601 ^ x239 ;
  assign n8603 = x535 ^ x240 ;
  assign n8604 = ~n6542 & n8603 ;
  assign n8605 = n8604 ^ x240 ;
  assign n8606 = x536 ^ x246 ;
  assign n8607 = ~n6542 & n8606 ;
  assign n8608 = n8607 ^ x246 ;
  assign n8609 = x537 ^ x248 ;
  assign n8610 = ~n6542 & n8609 ;
  assign n8611 = n8610 ^ x248 ;
  assign n8612 = x538 ^ x249 ;
  assign n8613 = ~n6542 & n8612 ;
  assign n8614 = n8613 ^ x249 ;
  assign n8615 = x539 ^ x242 ;
  assign n8616 = ~n6541 & n8615 ;
  assign n8617 = n8616 ^ x242 ;
  assign n8618 = x540 ^ x235 ;
  assign n8619 = ~n6541 & n8618 ;
  assign n8620 = n8619 ^ x235 ;
  assign n8621 = x541 ^ x244 ;
  assign n8622 = ~n6541 & n8621 ;
  assign n8623 = n8622 ^ x244 ;
  assign n8624 = x542 ^ x240 ;
  assign n8625 = ~n6541 & n8624 ;
  assign n8626 = n8625 ^ x240 ;
  assign n8627 = x543 ^ x238 ;
  assign n8628 = ~n6541 & n8627 ;
  assign n8629 = n8628 ^ x238 ;
  assign n8630 = x544 ^ x234 ;
  assign n8631 = ~n6556 & n8630 ;
  assign n8632 = n8631 ^ x234 ;
  assign n8633 = x545 ^ x245 ;
  assign n8634 = ~n6556 & n8633 ;
  assign n8635 = n8634 ^ x245 ;
  assign n8636 = x546 ^ x246 ;
  assign n8637 = ~n6556 & n8636 ;
  assign n8638 = n8637 ^ x246 ;
  assign n8639 = x547 ^ x247 ;
  assign n8640 = ~n6556 & n8639 ;
  assign n8641 = n8640 ^ x247 ;
  assign n8642 = x548 ^ x248 ;
  assign n8643 = ~n6556 & n8642 ;
  assign n8644 = n8643 ^ x248 ;
  assign n8645 = x549 ^ x235 ;
  assign n8646 = ~n6555 & n8645 ;
  assign n8647 = n8646 ^ x235 ;
  assign n8648 = x550 ^ x239 ;
  assign n8649 = ~n6555 & ~n8648 ;
  assign n8650 = n8649 ^ x239 ;
  assign n8651 = x551 ^ x240 ;
  assign n8652 = ~n6555 & n8651 ;
  assign n8653 = n8652 ^ x240 ;
  assign n8654 = x552 ^ x247 ;
  assign n8655 = ~n6555 & n8654 ;
  assign n8656 = n8655 ^ x247 ;
  assign n8657 = x553 ^ x241 ;
  assign n8658 = ~n6555 & n8657 ;
  assign n8659 = n8658 ^ x241 ;
  assign n8660 = x554 ^ x248 ;
  assign n8661 = ~n6555 & n8660 ;
  assign n8662 = n8661 ^ x248 ;
  assign n8663 = x555 ^ x249 ;
  assign n8664 = ~n6555 & n8663 ;
  assign n8665 = n8664 ^ x249 ;
  assign n8666 = x556 ^ x242 ;
  assign n8667 = ~n6524 & n8666 ;
  assign n8668 = n8667 ^ x242 ;
  assign n8669 = x557 ^ x234 ;
  assign n8670 = ~n6542 & n8669 ;
  assign n8671 = n8670 ^ x234 ;
  assign n8672 = x558 ^ x244 ;
  assign n8673 = ~n6542 & n8672 ;
  assign n8674 = n8673 ^ x244 ;
  assign n8675 = x559 ^ x241 ;
  assign n8676 = ~n6508 & n8675 ;
  assign n8677 = n8676 ^ x241 ;
  assign n8678 = x560 ^ x240 ;
  assign n8679 = ~n6524 & n8678 ;
  assign n8680 = n8679 ^ x240 ;
  assign n8681 = x561 ^ x247 ;
  assign n8682 = ~n6517 & n8681 ;
  assign n8683 = n8682 ^ x247 ;
  assign n8684 = x562 ^ x241 ;
  assign n8685 = ~n6524 & n8684 ;
  assign n8686 = n8685 ^ x241 ;
  assign n8687 = x563 ^ x246 ;
  assign n8688 = ~n6555 & n8687 ;
  assign n8689 = n8688 ^ x246 ;
  assign n8690 = x564 ^ x246 ;
  assign n8691 = ~n6524 & n8690 ;
  assign n8692 = n8691 ^ x246 ;
  assign n8693 = x565 ^ x248 ;
  assign n8694 = ~n6524 & n8693 ;
  assign n8695 = n8694 ^ x248 ;
  assign n8696 = x566 ^ x244 ;
  assign n8697 = ~n6524 & n8696 ;
  assign n8698 = n8697 ^ x244 ;
  assign n8699 = x230 & x1093 ;
  assign n8703 = n5837 ^ x567 ;
  assign n8700 = n5837 ^ x1091 ;
  assign n8701 = x621 & n5800 ;
  assign n8702 = n8700 & n8701 ;
  assign n8704 = n8703 ^ n8702 ;
  assign n8705 = n8699 & ~n8704 ;
  assign n8706 = n8705 ^ x567 ;
  assign n8707 = x1092 & ~n8706 ;
  assign n8708 = x568 ^ x245 ;
  assign n8709 = ~n6524 & n8708 ;
  assign n8710 = n8709 ^ x245 ;
  assign n8711 = x569 ^ x239 ;
  assign n8712 = ~n6524 & ~n8711 ;
  assign n8713 = n8712 ^ x239 ;
  assign n8714 = x570 ^ x234 ;
  assign n8715 = ~n6524 & n8714 ;
  assign n8716 = n8715 ^ x234 ;
  assign n8717 = x571 ^ x241 ;
  assign n8718 = ~n6690 & n8717 ;
  assign n8719 = n8718 ^ x241 ;
  assign n8720 = x572 ^ x244 ;
  assign n8721 = ~n6690 & n8720 ;
  assign n8722 = n8721 ^ x244 ;
  assign n8723 = x573 ^ x242 ;
  assign n8724 = ~n6690 & n8723 ;
  assign n8725 = n8724 ^ x242 ;
  assign n8726 = x574 ^ x241 ;
  assign n8727 = ~n6517 & n8726 ;
  assign n8728 = n8727 ^ x241 ;
  assign n8729 = x575 ^ x235 ;
  assign n8730 = ~n6690 & n8729 ;
  assign n8731 = n8730 ^ x235 ;
  assign n8732 = x576 ^ x248 ;
  assign n8733 = ~n6690 & n8732 ;
  assign n8734 = n8733 ^ x248 ;
  assign n8735 = x577 ^ x238 ;
  assign n8736 = ~n6555 & n8735 ;
  assign n8737 = n8736 ^ x238 ;
  assign n8738 = x578 ^ x249 ;
  assign n8739 = ~n6517 & n8738 ;
  assign n8740 = n8739 ^ x249 ;
  assign n8741 = x579 ^ x249 ;
  assign n8742 = ~n6508 & n8741 ;
  assign n8743 = n8742 ^ x249 ;
  assign n8744 = x580 ^ x245 ;
  assign n8745 = ~n6555 & n8744 ;
  assign n8746 = n8745 ^ x245 ;
  assign n8747 = x581 ^ x235 ;
  assign n8748 = ~n6517 & n8747 ;
  assign n8749 = n8748 ^ x235 ;
  assign n8750 = x582 ^ x240 ;
  assign n8751 = ~n6517 & n8750 ;
  assign n8752 = n8751 ^ x240 ;
  assign n8753 = x584 ^ x245 ;
  assign n8754 = ~n6517 & n8753 ;
  assign n8755 = n8754 ^ x245 ;
  assign n8756 = x585 ^ x244 ;
  assign n8757 = ~n6517 & n8756 ;
  assign n8758 = n8757 ^ x244 ;
  assign n8759 = x586 ^ x242 ;
  assign n8760 = ~n6517 & n8759 ;
  assign n8761 = n8760 ^ x242 ;
  assign n8762 = n5802 ^ x587 ;
  assign n8763 = x230 & n8762 ;
  assign n8764 = n8763 ^ x587 ;
  assign n8765 = x591 ^ x588 ;
  assign n8766 = ~x123 & x824 ;
  assign n8767 = x950 & n8766 ;
  assign n8770 = n8765 & ~n8767 ;
  assign n8771 = n8770 ^ x591 ;
  assign n8772 = n7929 & n8771 ;
  assign n8773 = x218 ^ x205 ;
  assign n8774 = ~x237 & n8773 ;
  assign n8775 = n8774 ^ x205 ;
  assign n8777 = n8775 ^ x204 ;
  assign n8776 = n8775 ^ x206 ;
  assign n8778 = n8777 ^ n8776 ;
  assign n8781 = x237 & n8778 ;
  assign n8782 = n8781 ^ n8776 ;
  assign n8783 = x233 & n8782 ;
  assign n8784 = n8783 ^ n8775 ;
  assign n8785 = n6538 & ~n8784 ;
  assign n8786 = x203 ^ x202 ;
  assign n8787 = ~x237 & n8786 ;
  assign n8788 = n8787 ^ x202 ;
  assign n8790 = n8788 ^ x201 ;
  assign n8789 = n8788 ^ x220 ;
  assign n8791 = n8790 ^ n8789 ;
  assign n8794 = x237 & n8791 ;
  assign n8795 = n8794 ^ n8789 ;
  assign n8796 = x233 & n8795 ;
  assign n8797 = n8796 ^ n8788 ;
  assign n8798 = n6501 & ~n8797 ;
  assign n8799 = ~n8785 & ~n8798 ;
  assign n8800 = x590 ^ x588 ;
  assign n8803 = n8767 & n8800 ;
  assign n8804 = n8803 ^ x590 ;
  assign n8805 = n7929 & ~n8804 ;
  assign n8806 = x592 ^ x591 ;
  assign n8809 = n8767 & n8806 ;
  assign n8810 = n8809 ^ x591 ;
  assign n8811 = n7929 & n8810 ;
  assign n8814 = n3078 & ~n8767 ;
  assign n8815 = n8814 ^ x590 ;
  assign n8816 = n7929 & n8815 ;
  assign n8844 = ~n8453 & ~n8687 ;
  assign n8845 = ~n8735 & ~n8744 ;
  assign n8846 = n8844 & n8845 ;
  assign n8847 = ~n8645 & n8648 ;
  assign n8848 = ~n8657 & ~n8663 ;
  assign n8849 = n8847 & n8848 ;
  assign n8850 = n8846 & n8849 ;
  assign n8851 = ~n8456 & ~n8651 ;
  assign n8852 = ~x233 & ~n8465 ;
  assign n8853 = ~n8654 & ~n8660 ;
  assign n8854 = n8852 & n8853 ;
  assign n8855 = n8851 & n8854 ;
  assign n8856 = n8850 & n8855 ;
  assign n8857 = ~n8450 & ~n8477 ;
  assign n8858 = ~n8636 & ~n8642 ;
  assign n8859 = n8857 & n8858 ;
  assign n8860 = ~n8474 & n8480 ;
  assign n8861 = ~n8483 & ~n8630 ;
  assign n8862 = n8860 & n8861 ;
  assign n8863 = n8859 & n8862 ;
  assign n8864 = ~n8447 & ~n8471 ;
  assign n8865 = x233 & ~n8468 ;
  assign n8866 = ~n8633 & ~n8639 ;
  assign n8867 = n8865 & n8866 ;
  assign n8868 = n8864 & n8867 ;
  assign n8869 = n8863 & n8868 ;
  assign n8870 = ~n8856 & ~n8869 ;
  assign n8817 = ~n8516 & ~n8603 ;
  assign n8818 = ~n8669 & ~n8672 ;
  assign n8819 = n8817 & n8818 ;
  assign n8820 = ~n8525 & n8600 ;
  assign n8821 = ~n8606 & ~n8609 ;
  assign n8822 = n8820 & n8821 ;
  assign n8823 = n8819 & n8822 ;
  assign n8824 = ~n8510 & ~n8522 ;
  assign n8825 = x233 & ~n8519 ;
  assign n8826 = ~n8597 & ~n8612 ;
  assign n8827 = n8825 & n8826 ;
  assign n8828 = n8824 & n8827 ;
  assign n8829 = n8823 & n8828 ;
  assign n8830 = ~n8501 & ~n8504 ;
  assign n8831 = ~n8618 & ~n8627 ;
  assign n8832 = n8830 & n8831 ;
  assign n8833 = n8489 & ~n8513 ;
  assign n8834 = ~n8621 & ~n8624 ;
  assign n8835 = n8833 & n8834 ;
  assign n8836 = n8832 & n8835 ;
  assign n8837 = ~n8507 & ~n8615 ;
  assign n8838 = ~x233 & ~n8486 ;
  assign n8839 = ~n8498 & n8838 ;
  assign n8840 = n8837 & n8839 ;
  assign n8841 = ~n8495 & n8840 ;
  assign n8842 = n8836 & n8841 ;
  assign n8843 = ~n8829 & ~n8842 ;
  assign n8871 = n8870 ^ n8843 ;
  assign n8872 = x237 & n8871 ;
  assign n8873 = n8872 ^ n8870 ;
  assign n8874 = n6538 & ~n8873 ;
  assign n8902 = n8570 & ~n8573 ;
  assign n8903 = ~n8582 & ~n8585 ;
  assign n8904 = n8902 & n8903 ;
  assign n8905 = ~n8567 & ~n8576 ;
  assign n8906 = ~n8723 & ~n8729 ;
  assign n8907 = n8905 & n8906 ;
  assign n8908 = n8904 & n8907 ;
  assign n8909 = x233 & ~n8717 ;
  assign n8910 = x244 & ~x572 ;
  assign n8911 = n8910 ^ n8720 ;
  assign n8912 = ~n8579 & ~n8732 ;
  assign n8913 = ~n8911 & n8912 ;
  assign n8914 = n8909 & n8913 ;
  assign n8915 = n8908 & n8914 ;
  assign n8916 = ~n8588 & ~n8910 ;
  assign n8917 = n8915 & n8916 ;
  assign n8918 = ~n8693 & ~n8714 ;
  assign n8919 = ~n8678 & ~n8690 ;
  assign n8920 = n8918 & n8919 ;
  assign n8921 = ~n8492 & ~n8594 ;
  assign n8922 = ~n8708 & n8711 ;
  assign n8923 = n8921 & n8922 ;
  assign n8924 = n8920 & n8923 ;
  assign n8925 = ~n8591 & ~n8696 ;
  assign n8926 = x249 & ~x482 ;
  assign n8927 = n8926 ^ n8444 ;
  assign n8928 = ~x233 & ~n8684 ;
  assign n8929 = ~n8927 & n8928 ;
  assign n8930 = n8925 & n8929 ;
  assign n8931 = n8924 & n8930 ;
  assign n8932 = ~n8666 & ~n8926 ;
  assign n8933 = n8931 & n8932 ;
  assign n8934 = ~n8917 & ~n8933 ;
  assign n8875 = ~n8528 & ~n8531 ;
  assign n8876 = ~n8537 & ~n8543 ;
  assign n8877 = n8875 & n8876 ;
  assign n8878 = ~n8459 & n8462 ;
  assign n8879 = ~n8534 & ~n8549 ;
  assign n8880 = n8878 & n8879 ;
  assign n8881 = n8877 & n8880 ;
  assign n8882 = ~n8441 & ~n8546 ;
  assign n8883 = x233 & ~n8540 ;
  assign n8884 = ~n8675 & ~n8741 ;
  assign n8885 = n8883 & n8884 ;
  assign n8886 = n8882 & n8885 ;
  assign n8887 = n8881 & n8886 ;
  assign n8888 = ~n8552 & n8555 ;
  assign n8889 = ~n8558 & ~n8753 ;
  assign n8890 = n8888 & n8889 ;
  assign n8891 = ~n8681 & ~n8747 ;
  assign n8892 = ~n8750 & ~n8759 ;
  assign n8893 = n8891 & n8892 ;
  assign n8894 = n8890 & n8893 ;
  assign n8895 = ~n8561 & ~n8726 ;
  assign n8896 = ~x233 & ~n8564 ;
  assign n8897 = ~n8738 & ~n8756 ;
  assign n8898 = n8896 & n8897 ;
  assign n8899 = n8895 & n8898 ;
  assign n8900 = n8894 & n8899 ;
  assign n8901 = ~n8887 & ~n8900 ;
  assign n8935 = n8934 ^ n8901 ;
  assign n8936 = x237 & n8935 ;
  assign n8937 = n8936 ^ n8934 ;
  assign n8938 = n6501 & ~n8937 ;
  assign n8939 = ~n8874 & ~n8938 ;
  assign n8940 = ~x806 & x990 ;
  assign n8945 = x600 & n8940 ;
  assign n8946 = n8945 ^ x594 ;
  assign n8947 = ~x332 & n8946 ;
  assign n8954 = ~x806 & n8316 ;
  assign n8955 = x605 & n8954 ;
  assign n8956 = n8955 ^ x605 ;
  assign n8948 = x605 ^ x595 ;
  assign n8957 = n8956 ^ n8948 ;
  assign n8958 = ~x332 & n8957 ;
  assign n8959 = n8314 & n8940 ;
  assign n8960 = x595 & x597 ;
  assign n8961 = n8959 & n8960 ;
  assign n8962 = n8961 ^ x596 ;
  assign n8963 = ~x332 & n8962 ;
  assign n8964 = n8959 ^ x597 ;
  assign n8965 = ~x332 & n8964 ;
  assign n8966 = ~x882 & n1290 ;
  assign n8967 = x947 & n8966 ;
  assign n8968 = x598 & ~n8967 ;
  assign n8969 = x740 & x780 ;
  assign n8970 = n2665 & n8969 ;
  assign n8971 = n8968 & ~n8970 ;
  assign n8972 = n8971 ^ n8970 ;
  assign n8977 = x596 & n8961 ;
  assign n8978 = n8977 ^ x599 ;
  assign n8979 = ~x332 & n8978 ;
  assign n8980 = n8940 ^ x600 ;
  assign n8981 = ~x332 & n8980 ;
  assign n8982 = x989 ^ x601 ;
  assign n8983 = ~x806 & n8982 ;
  assign n8984 = n8983 ^ x601 ;
  assign n8985 = ~x332 & n8984 ;
  assign n8986 = n5838 ^ x602 ;
  assign n8987 = x230 & n8986 ;
  assign n8988 = n8987 ^ x602 ;
  assign n9002 = ~x871 & ~x872 ;
  assign n8989 = x1100 ^ x603 ;
  assign n8990 = x832 & ~x980 ;
  assign n8991 = x1060 & n8990 ;
  assign n8992 = x1038 & ~x1061 ;
  assign n8993 = n8991 & n8992 ;
  assign n8994 = ~x952 & n8993 ;
  assign n8995 = n8994 ^ n8993 ;
  assign n8996 = n8989 & n8995 ;
  assign n8997 = n8996 ^ x603 ;
  assign n9003 = n9002 ^ n8997 ;
  assign n9004 = x966 & ~n9003 ;
  assign n9005 = n9004 ^ n8997 ;
  assign n9006 = x823 & n2667 ;
  assign n9010 = ~x299 & x983 ;
  assign n9015 = x604 & n9010 ;
  assign n9016 = x907 & n9015 ;
  assign n9017 = n9016 ^ x907 ;
  assign n9007 = x779 ^ x604 ;
  assign n9008 = n9007 ^ x907 ;
  assign n9018 = n9017 ^ n9008 ;
  assign n9019 = ~n9006 & ~n9018 ;
  assign n9020 = n9019 ^ x779 ;
  assign n9021 = x806 ^ x605 ;
  assign n9022 = ~x332 & ~n9021 ;
  assign n9026 = x1104 ^ x837 ;
  assign n9023 = x837 ^ x606 ;
  assign n9027 = n9026 ^ n9023 ;
  assign n9028 = n8995 & n9027 ;
  assign n9029 = n9028 ^ n9023 ;
  assign n9030 = ~x966 & n9029 ;
  assign n9031 = n9030 ^ x837 ;
  assign n9032 = x1107 ^ x607 ;
  assign n9035 = n8995 & n9032 ;
  assign n9036 = n9035 ^ x607 ;
  assign n9037 = ~x966 & n9036 ;
  assign n9038 = x1116 ^ x608 ;
  assign n9041 = n8995 & n9038 ;
  assign n9042 = n9041 ^ x608 ;
  assign n9043 = ~x966 & n9042 ;
  assign n9044 = x1118 ^ x609 ;
  assign n9047 = n8995 & n9044 ;
  assign n9048 = n9047 ^ x609 ;
  assign n9049 = ~x966 & n9048 ;
  assign n9050 = x1113 ^ x610 ;
  assign n9053 = n8995 & n9050 ;
  assign n9054 = n9053 ^ x610 ;
  assign n9055 = ~x966 & n9054 ;
  assign n9056 = x1114 ^ x611 ;
  assign n9059 = n8995 & n9056 ;
  assign n9060 = n9059 ^ x611 ;
  assign n9061 = ~x966 & n9060 ;
  assign n9062 = x1111 ^ x612 ;
  assign n9065 = n8995 & n9062 ;
  assign n9066 = n9065 ^ x612 ;
  assign n9067 = ~x966 & n9066 ;
  assign n9068 = x1115 ^ x613 ;
  assign n9071 = n8995 & n9068 ;
  assign n9072 = n9071 ^ x613 ;
  assign n9073 = ~x966 & n9072 ;
  assign n9077 = x1102 ^ x871 ;
  assign n9074 = x871 ^ x614 ;
  assign n9078 = n9077 ^ n9074 ;
  assign n9079 = n8995 & n9078 ;
  assign n9080 = n9079 ^ n9074 ;
  assign n9081 = ~x966 & n9080 ;
  assign n9082 = n9081 ^ x871 ;
  assign n9083 = x907 & n8966 ;
  assign n9084 = ~x615 & ~n9083 ;
  assign n9085 = x779 & x797 ;
  assign n9086 = n2668 & n9085 ;
  assign n9087 = n9084 & ~n9086 ;
  assign n9088 = n9087 ^ n9086 ;
  assign n9092 = x1101 ^ x872 ;
  assign n9089 = x872 ^ x616 ;
  assign n9093 = n9092 ^ n9089 ;
  assign n9094 = n8995 & n9093 ;
  assign n9095 = n9094 ^ n9089 ;
  assign n9096 = ~x966 & n9095 ;
  assign n9097 = n9096 ^ x872 ;
  assign n9101 = x1105 ^ x850 ;
  assign n9098 = x850 ^ x617 ;
  assign n9102 = n9101 ^ n9098 ;
  assign n9103 = n8995 & n9102 ;
  assign n9104 = n9103 ^ n9098 ;
  assign n9105 = ~x966 & n9104 ;
  assign n9106 = n9105 ^ x850 ;
  assign n9107 = x1117 ^ x618 ;
  assign n9110 = n8995 & n9107 ;
  assign n9111 = n9110 ^ x618 ;
  assign n9112 = ~x966 & n9111 ;
  assign n9113 = x1122 ^ x619 ;
  assign n9116 = n8995 & n9113 ;
  assign n9117 = n9116 ^ x619 ;
  assign n9118 = ~x966 & n9117 ;
  assign n9119 = x1112 ^ x620 ;
  assign n9122 = n8995 & n9119 ;
  assign n9123 = n9122 ^ x620 ;
  assign n9124 = ~x966 & n9123 ;
  assign n9125 = x1108 ^ x621 ;
  assign n9128 = n8995 & n9125 ;
  assign n9129 = n9128 ^ x621 ;
  assign n9130 = ~x966 & n9129 ;
  assign n9131 = x1109 ^ x622 ;
  assign n9134 = n8995 & n9131 ;
  assign n9135 = n9134 ^ x622 ;
  assign n9136 = ~x966 & n9135 ;
  assign n9137 = x1106 ^ x623 ;
  assign n9140 = n8995 & n9137 ;
  assign n9141 = n9140 ^ x623 ;
  assign n9142 = ~x966 & n9141 ;
  assign n9143 = x831 & n2664 ;
  assign n9151 = x624 & n9010 ;
  assign n9152 = x947 & n9151 ;
  assign n9153 = n9152 ^ x947 ;
  assign n9144 = x780 ^ x624 ;
  assign n9145 = n9144 ^ x947 ;
  assign n9154 = n9153 ^ n9145 ;
  assign n9155 = ~n9143 & ~n9154 ;
  assign n9156 = n9155 ^ x780 ;
  assign n9157 = x1116 ^ x625 ;
  assign n9158 = x1066 & x1088 ;
  assign n9159 = ~x973 & ~x1054 ;
  assign n9160 = n9158 & n9159 ;
  assign n9161 = x832 & n9160 ;
  assign n9162 = x953 & n9161 ;
  assign n9163 = n9162 ^ n9161 ;
  assign n9166 = n9157 & n9163 ;
  assign n9167 = n9166 ^ x625 ;
  assign n9168 = ~x962 & n9167 ;
  assign n9169 = x1121 ^ x626 ;
  assign n9172 = n8995 & n9169 ;
  assign n9173 = n9172 ^ x626 ;
  assign n9174 = ~x966 & n9173 ;
  assign n9175 = x1117 ^ x627 ;
  assign n9178 = n9163 & n9175 ;
  assign n9179 = n9178 ^ x627 ;
  assign n9180 = ~x962 & n9179 ;
  assign n9181 = x1119 ^ x628 ;
  assign n9184 = n9163 & n9181 ;
  assign n9185 = n9184 ^ x628 ;
  assign n9186 = ~x962 & n9185 ;
  assign n9187 = x1119 ^ x629 ;
  assign n9190 = n8995 & n9187 ;
  assign n9191 = n9190 ^ x629 ;
  assign n9192 = ~x966 & n9191 ;
  assign n9193 = x1120 ^ x630 ;
  assign n9196 = n8995 & n9193 ;
  assign n9197 = n9196 ^ x630 ;
  assign n9198 = ~x966 & n9197 ;
  assign n9199 = x1113 ^ x631 ;
  assign n9202 = n9163 & ~n9199 ;
  assign n9203 = n9202 ^ x631 ;
  assign n9204 = ~x962 & ~n9203 ;
  assign n9205 = x1115 ^ x632 ;
  assign n9208 = n9163 & ~n9205 ;
  assign n9209 = n9208 ^ x632 ;
  assign n9210 = ~x962 & ~n9209 ;
  assign n9211 = x1110 ^ x633 ;
  assign n9214 = n8995 & n9211 ;
  assign n9215 = n9214 ^ x633 ;
  assign n9216 = ~x966 & n9215 ;
  assign n9217 = x1110 ^ x634 ;
  assign n9220 = n9163 & n9217 ;
  assign n9221 = n9220 ^ x634 ;
  assign n9222 = ~x962 & n9221 ;
  assign n9223 = x1112 ^ x635 ;
  assign n9226 = n9163 & ~n9223 ;
  assign n9227 = n9226 ^ x635 ;
  assign n9228 = ~x962 & ~n9227 ;
  assign n9229 = x1127 ^ x636 ;
  assign n9232 = n8995 & n9229 ;
  assign n9233 = n9232 ^ x636 ;
  assign n9234 = ~x966 & n9233 ;
  assign n9235 = x1105 ^ x637 ;
  assign n9238 = n9163 & n9235 ;
  assign n9239 = n9238 ^ x637 ;
  assign n9240 = ~x962 & n9239 ;
  assign n9241 = x1107 ^ x638 ;
  assign n9244 = n9163 & n9241 ;
  assign n9245 = n9244 ^ x638 ;
  assign n9246 = ~x962 & n9245 ;
  assign n9247 = x1109 ^ x639 ;
  assign n9250 = n9163 & n9247 ;
  assign n9251 = n9250 ^ x639 ;
  assign n9252 = ~x962 & n9251 ;
  assign n9253 = x1128 ^ x640 ;
  assign n9256 = n8995 & n9253 ;
  assign n9257 = n9256 ^ x640 ;
  assign n9258 = ~x966 & n9257 ;
  assign n9259 = x1121 ^ x641 ;
  assign n9262 = n9163 & n9259 ;
  assign n9263 = n9262 ^ x641 ;
  assign n9264 = ~x962 & n9263 ;
  assign n9265 = x1103 ^ x642 ;
  assign n9268 = n8995 & n9265 ;
  assign n9269 = n9268 ^ x642 ;
  assign n9270 = ~x966 & n9269 ;
  assign n9271 = x1104 ^ x643 ;
  assign n9274 = n9163 & n9271 ;
  assign n9275 = n9274 ^ x643 ;
  assign n9276 = ~x962 & n9275 ;
  assign n9277 = x1123 ^ x644 ;
  assign n9280 = n8995 & n9277 ;
  assign n9281 = n9280 ^ x644 ;
  assign n9282 = ~x966 & n9281 ;
  assign n9283 = x1125 ^ x645 ;
  assign n9286 = n8995 & n9283 ;
  assign n9287 = n9286 ^ x645 ;
  assign n9288 = ~x966 & n9287 ;
  assign n9289 = x1114 ^ x646 ;
  assign n9292 = n9163 & ~n9289 ;
  assign n9293 = n9292 ^ x646 ;
  assign n9294 = ~x962 & ~n9293 ;
  assign n9295 = x1120 ^ x647 ;
  assign n9298 = n9163 & n9295 ;
  assign n9299 = n9298 ^ x647 ;
  assign n9300 = ~x962 & n9299 ;
  assign n9301 = x1122 ^ x648 ;
  assign n9304 = n9163 & n9301 ;
  assign n9305 = n9304 ^ x648 ;
  assign n9306 = ~x962 & n9305 ;
  assign n9307 = x1126 ^ x649 ;
  assign n9310 = n9163 & ~n9307 ;
  assign n9311 = n9310 ^ x649 ;
  assign n9312 = ~x962 & ~n9311 ;
  assign n9313 = x1127 ^ x650 ;
  assign n9316 = n9163 & ~n9313 ;
  assign n9317 = n9316 ^ x650 ;
  assign n9318 = ~x962 & ~n9317 ;
  assign n9319 = x1130 ^ x651 ;
  assign n9322 = n8995 & n9319 ;
  assign n9323 = n9322 ^ x651 ;
  assign n9324 = ~x966 & n9323 ;
  assign n9325 = x1131 ^ x652 ;
  assign n9328 = n8995 & n9325 ;
  assign n9329 = n9328 ^ x652 ;
  assign n9330 = ~x966 & n9329 ;
  assign n9331 = x1129 ^ x653 ;
  assign n9334 = n8995 & n9331 ;
  assign n9335 = n9334 ^ x653 ;
  assign n9336 = ~x966 & n9335 ;
  assign n9337 = x1130 ^ x654 ;
  assign n9340 = n9163 & ~n9337 ;
  assign n9341 = n9340 ^ x654 ;
  assign n9342 = ~x962 & ~n9341 ;
  assign n9343 = x1124 ^ x655 ;
  assign n9346 = n9163 & ~n9343 ;
  assign n9347 = n9346 ^ x655 ;
  assign n9348 = ~x962 & ~n9347 ;
  assign n9349 = x1126 ^ x656 ;
  assign n9352 = n8995 & n9349 ;
  assign n9353 = n9352 ^ x656 ;
  assign n9354 = ~x966 & n9353 ;
  assign n9355 = x1131 ^ x657 ;
  assign n9358 = n9163 & ~n9355 ;
  assign n9359 = n9358 ^ x657 ;
  assign n9360 = ~x962 & ~n9359 ;
  assign n9361 = x1124 ^ x658 ;
  assign n9364 = n8995 & n9361 ;
  assign n9365 = n9364 ^ x658 ;
  assign n9366 = ~x966 & n9365 ;
  assign n9367 = x266 & x992 ;
  assign n9368 = ~x280 & n9367 ;
  assign n9369 = ~x269 & n9368 ;
  assign n9370 = ~x281 & ~x282 ;
  assign n9371 = n9369 & n9370 ;
  assign n9372 = ~x270 & ~x277 ;
  assign n9373 = ~x264 & n9372 ;
  assign n9374 = n9371 & n9373 ;
  assign n9375 = ~x265 & n9374 ;
  assign n9376 = n9375 ^ x274 ;
  assign n9377 = x1118 ^ x660 ;
  assign n9380 = n9163 & n9377 ;
  assign n9381 = n9380 ^ x660 ;
  assign n9382 = ~x962 & n9381 ;
  assign n9383 = x1101 ^ x661 ;
  assign n9386 = n9163 & n9383 ;
  assign n9387 = n9386 ^ x661 ;
  assign n9388 = ~x962 & n9387 ;
  assign n9389 = x1102 ^ x662 ;
  assign n9392 = n9163 & n9389 ;
  assign n9393 = n9392 ^ x662 ;
  assign n9394 = ~x962 & n9393 ;
  assign n9395 = ~x1137 & ~x1138 ;
  assign n9396 = ~n3209 & n9395 ;
  assign n9406 = x815 ^ x633 ;
  assign n9407 = ~x1136 & n9406 ;
  assign n9408 = n9407 ^ x633 ;
  assign n9410 = n9408 ^ x766 ;
  assign n9409 = n9408 ^ x855 ;
  assign n9411 = n9410 ^ n9409 ;
  assign n9414 = x1136 & n9411 ;
  assign n9415 = n9414 ^ n9409 ;
  assign n9416 = x1134 & n9415 ;
  assign n9417 = n9416 ^ n9408 ;
  assign n9398 = x1135 ^ x1134 ;
  assign n9399 = x700 ^ x634 ;
  assign n9400 = n9399 ^ x784 ;
  assign n9403 = x1136 & n9400 ;
  assign n9404 = n9403 ^ x784 ;
  assign n9405 = n9398 & n9404 ;
  assign n9418 = n9417 ^ n9405 ;
  assign n9397 = x700 & x1136 ;
  assign n9419 = n9418 ^ n9397 ;
  assign n9420 = x1135 & n9419 ;
  assign n9421 = n9420 ^ n9417 ;
  assign n9422 = n9396 & n9421 ;
  assign n9423 = ~x223 & ~x224 ;
  assign n9424 = n4592 & n8806 ;
  assign n9425 = n9423 & n9424 ;
  assign n9426 = x365 ^ x334 ;
  assign n9429 = ~x592 & n9426 ;
  assign n9430 = n9429 ^ x365 ;
  assign n9431 = n9425 & n9430 ;
  assign n9432 = n9431 ^ n9423 ;
  assign n9433 = ~x591 & n3015 ;
  assign n9435 = ~x588 & ~n9433 ;
  assign n9434 = n9433 ^ x588 ;
  assign n9436 = n9435 ^ n9434 ;
  assign n9437 = x464 & ~n9436 ;
  assign n9438 = n9432 & n9437 ;
  assign n9439 = n9438 ^ x323 ;
  assign n9441 = n9435 & n9440 ;
  assign n9442 = n9438 ^ n9432 ;
  assign n9443 = n3209 & ~n9423 ;
  assign n9444 = x1065 ^ x257 ;
  assign n9447 = x199 & n9444 ;
  assign n9448 = n9447 ^ x257 ;
  assign n9449 = n9443 & ~n9448 ;
  assign n9450 = n9449 ^ n3209 ;
  assign n9451 = n9442 & n9450 ;
  assign n9452 = n9441 & n9451 ;
  assign n9453 = n9439 & n9452 ;
  assign n9454 = n9453 ^ n9451 ;
  assign n9455 = n9454 ^ n9450 ;
  assign n9456 = ~n9422 & ~n9455 ;
  assign n9465 = x811 ^ x614 ;
  assign n9466 = ~x1136 & n9465 ;
  assign n9467 = n9466 ^ x614 ;
  assign n9469 = n9467 ^ x772 ;
  assign n9468 = n9467 ^ x872 ;
  assign n9470 = n9469 ^ n9468 ;
  assign n9473 = x1136 & n9470 ;
  assign n9474 = n9473 ^ n9468 ;
  assign n9475 = x1134 & n9474 ;
  assign n9476 = n9475 ^ n9467 ;
  assign n9458 = x727 ^ x662 ;
  assign n9459 = n9458 ^ x785 ;
  assign n9462 = x1136 & n9459 ;
  assign n9463 = n9462 ^ x785 ;
  assign n9464 = n9398 & n9463 ;
  assign n9477 = n9476 ^ n9464 ;
  assign n9457 = x727 & x1136 ;
  assign n9478 = n9477 ^ n9457 ;
  assign n9479 = x1135 & n9478 ;
  assign n9480 = n9479 ^ n9476 ;
  assign n9481 = n9396 & n9480 ;
  assign n9488 = x404 ^ x380 ;
  assign n9491 = x592 & n9488 ;
  assign n9492 = n9491 ^ x404 ;
  assign n9493 = n9425 & n9492 ;
  assign n9494 = n9493 ^ n9423 ;
  assign n9495 = x429 & ~n9436 ;
  assign n9496 = n9494 & n9495 ;
  assign n9497 = n9496 ^ x355 ;
  assign n9484 = x199 & n7771 ;
  assign n9485 = n9484 ^ x292 ;
  assign n9486 = n9443 & ~n9485 ;
  assign n9487 = n9486 ^ n3209 ;
  assign n9498 = n9496 ^ n9494 ;
  assign n9499 = n9487 & n9498 ;
  assign n9500 = n9441 & n9499 ;
  assign n9501 = n9497 & n9500 ;
  assign n9502 = n9501 ^ n9499 ;
  assign n9503 = n9502 ^ n9487 ;
  assign n9504 = ~n9481 & ~n9503 ;
  assign n9505 = x1108 ^ x665 ;
  assign n9508 = n9163 & n9505 ;
  assign n9509 = n9508 ^ x665 ;
  assign n9510 = ~x962 & n9509 ;
  assign n9519 = x799 ^ x607 ;
  assign n9520 = ~x1136 & ~n9519 ;
  assign n9521 = n9520 ^ x607 ;
  assign n9523 = n9521 ^ x764 ;
  assign n9522 = n9521 ^ x873 ;
  assign n9524 = n9523 ^ n9522 ;
  assign n9527 = x1136 & n9524 ;
  assign n9528 = n9527 ^ n9522 ;
  assign n9529 = x1134 & n9528 ;
  assign n9530 = n9529 ^ n9521 ;
  assign n9512 = x691 ^ x638 ;
  assign n9513 = n9512 ^ x790 ;
  assign n9516 = x1136 & n9513 ;
  assign n9517 = n9516 ^ x790 ;
  assign n9518 = n9398 & n9517 ;
  assign n9531 = n9530 ^ n9518 ;
  assign n9511 = x691 & x1136 ;
  assign n9532 = n9531 ^ n9511 ;
  assign n9533 = x1135 & n9532 ;
  assign n9534 = n9533 ^ n9530 ;
  assign n9535 = n9396 & n9534 ;
  assign n9542 = x456 ^ x337 ;
  assign n9545 = x592 & n9542 ;
  assign n9546 = n9545 ^ x456 ;
  assign n9547 = n9425 & n9546 ;
  assign n9548 = n9547 ^ n9423 ;
  assign n9549 = x443 & ~n9436 ;
  assign n9550 = n9548 & n9549 ;
  assign n9551 = n9550 ^ x441 ;
  assign n9538 = x199 & n7786 ;
  assign n9539 = n9538 ^ x297 ;
  assign n9540 = n9443 & ~n9539 ;
  assign n9541 = n9540 ^ n3209 ;
  assign n9552 = n9550 ^ n9548 ;
  assign n9553 = n9541 & n9552 ;
  assign n9554 = n9441 & n9553 ;
  assign n9555 = n9551 & n9554 ;
  assign n9556 = n9555 ^ n9553 ;
  assign n9557 = n9556 ^ n9541 ;
  assign n9558 = ~n9535 & ~n9557 ;
  assign n9588 = x809 ^ x642 ;
  assign n9589 = ~x1136 & ~n9588 ;
  assign n9590 = n9589 ^ x642 ;
  assign n9592 = n9590 ^ x763 ;
  assign n9591 = n9590 ^ x871 ;
  assign n9593 = n9592 ^ n9591 ;
  assign n9596 = x1136 & n9593 ;
  assign n9597 = n9596 ^ n9591 ;
  assign n9598 = x1134 & n9597 ;
  assign n9599 = n9598 ^ n9590 ;
  assign n9581 = x699 ^ x681 ;
  assign n9582 = n9581 ^ x792 ;
  assign n9585 = x1136 & n9582 ;
  assign n9586 = n9585 ^ x792 ;
  assign n9587 = n9398 & n9586 ;
  assign n9600 = n9599 ^ n9587 ;
  assign n9580 = x699 & x1136 ;
  assign n9601 = n9600 ^ n9580 ;
  assign n9602 = x1135 & n9601 ;
  assign n9603 = n9602 ^ n9599 ;
  assign n9604 = n9395 & n9603 ;
  assign n9559 = x338 ^ x319 ;
  assign n9562 = ~x592 & n9559 ;
  assign n9563 = n9562 ^ x338 ;
  assign n9564 = n9424 & n9563 ;
  assign n9565 = n9564 ^ x444 ;
  assign n9570 = ~n9436 & n9565 ;
  assign n9566 = x458 & n9441 ;
  assign n9568 = n9566 ^ n9564 ;
  assign n9571 = n9570 ^ n9568 ;
  assign n9605 = n9604 ^ n9571 ;
  assign n9577 = x199 & n7777 ;
  assign n9573 = n9571 ^ x294 ;
  assign n9578 = n9577 ^ n9573 ;
  assign n9579 = ~n9423 & n9578 ;
  assign n9606 = n9605 ^ n9579 ;
  assign n9607 = n3209 & n9606 ;
  assign n9608 = n9607 ^ n9604 ;
  assign n9638 = x981 ^ x603 ;
  assign n9639 = ~x1136 & n9638 ;
  assign n9640 = n9639 ^ x603 ;
  assign n9642 = n9640 ^ x759 ;
  assign n9641 = n9640 ^ x837 ;
  assign n9643 = n9642 ^ n9641 ;
  assign n9646 = x1136 & n9643 ;
  assign n9647 = n9646 ^ n9641 ;
  assign n9648 = x1134 & n9647 ;
  assign n9649 = n9648 ^ n9640 ;
  assign n9631 = x696 ^ x680 ;
  assign n9632 = n9631 ^ x778 ;
  assign n9635 = x1136 & n9632 ;
  assign n9636 = n9635 ^ x778 ;
  assign n9637 = n9398 & n9636 ;
  assign n9650 = n9649 ^ n9637 ;
  assign n9630 = x696 & x1136 ;
  assign n9651 = n9650 ^ n9630 ;
  assign n9652 = x1135 & n9651 ;
  assign n9653 = n9652 ^ n9649 ;
  assign n9654 = n9395 & n9653 ;
  assign n9609 = x390 ^ x363 ;
  assign n9612 = x592 & n9609 ;
  assign n9613 = n9612 ^ x390 ;
  assign n9614 = n9424 & n9613 ;
  assign n9615 = n9614 ^ x342 ;
  assign n9620 = n9441 & n9615 ;
  assign n9616 = x414 & ~n9436 ;
  assign n9618 = n9616 ^ n9614 ;
  assign n9621 = n9620 ^ n9618 ;
  assign n9655 = n9654 ^ n9621 ;
  assign n9627 = x199 & n7768 ;
  assign n9623 = n9621 ^ x291 ;
  assign n9628 = n9627 ^ n9623 ;
  assign n9629 = ~n9423 & n9628 ;
  assign n9656 = n9655 ^ n9629 ;
  assign n9657 = n3209 & n9656 ;
  assign n9658 = n9657 ^ n9654 ;
  assign n9659 = x1125 ^ x669 ;
  assign n9662 = n9163 & ~n9659 ;
  assign n9663 = n9662 ^ x669 ;
  assign n9664 = ~x962 & ~n9663 ;
  assign n9678 = x1134 & ~x1135 ;
  assign n9679 = x852 & n9678 ;
  assign n5969 = x745 ^ x723 ;
  assign n9665 = ~x1135 & n5969 ;
  assign n9666 = n9665 ^ x723 ;
  assign n9668 = n9666 ^ x612 ;
  assign n9667 = n9666 ^ x695 ;
  assign n9669 = n9668 ^ n9667 ;
  assign n9672 = ~x1135 & ~n9669 ;
  assign n9673 = n9672 ^ n9667 ;
  assign n9674 = ~x1134 & n9673 ;
  assign n9675 = n9674 ^ n9666 ;
  assign n9680 = n9679 ^ n9675 ;
  assign n9681 = ~x1136 & ~n9680 ;
  assign n9682 = n9681 ^ n9675 ;
  assign n9683 = n9396 & ~n9682 ;
  assign n9684 = x1062 ^ x258 ;
  assign n9687 = x199 & n9684 ;
  assign n9688 = n9687 ^ x258 ;
  assign n9689 = n9443 & ~n9688 ;
  assign n9690 = n9689 ^ n3209 ;
  assign n9710 = x343 & n9441 ;
  assign n9711 = n9710 ^ x343 ;
  assign n9691 = x391 & ~x590 ;
  assign n9692 = ~x592 & n9691 ;
  assign n9693 = n9692 ^ x364 ;
  assign n9696 = n9692 ^ x590 ;
  assign n9697 = ~x591 & ~n9696 ;
  assign n9698 = n9693 & n9697 ;
  assign n9699 = n9698 ^ n9693 ;
  assign n9700 = n9699 ^ x364 ;
  assign n9701 = n9435 & ~n9700 ;
  assign n9702 = n9701 ^ n9435 ;
  assign n9703 = n9702 ^ x343 ;
  assign n9712 = n9711 ^ n9703 ;
  assign n9713 = n9423 & ~n9712 ;
  assign n9714 = n9690 & n9713 ;
  assign n9722 = x415 & n9714 ;
  assign n9723 = ~n9436 & n9722 ;
  assign n9724 = n9723 ^ n9436 ;
  assign n9715 = n9714 ^ n9690 ;
  assign n9716 = n9715 ^ n9436 ;
  assign n9725 = n9724 ^ n9716 ;
  assign n9726 = ~n9683 & ~n9725 ;
  assign n9727 = x447 ^ x333 ;
  assign n9730 = ~x592 & n9727 ;
  assign n9731 = n9730 ^ x447 ;
  assign n9732 = n9425 & n9731 ;
  assign n9733 = n9732 ^ n9423 ;
  assign n9734 = x453 & ~n9436 ;
  assign n9735 = n9733 & n9734 ;
  assign n9736 = n9735 ^ x327 ;
  assign n9737 = n9735 ^ n9733 ;
  assign n9738 = x1040 ^ x261 ;
  assign n9741 = x199 & n9738 ;
  assign n9742 = n9741 ^ x261 ;
  assign n9743 = n9443 & ~n9742 ;
  assign n9744 = n9743 ^ n3209 ;
  assign n9745 = n9737 & n9744 ;
  assign n9746 = n9441 & n9745 ;
  assign n9747 = n9736 & n9746 ;
  assign n9748 = n9747 ^ n9745 ;
  assign n9749 = n9748 ^ n9744 ;
  assign n9763 = x865 & n9678 ;
  assign n6028 = x741 ^ x724 ;
  assign n9750 = ~x1135 & n6028 ;
  assign n9751 = n9750 ^ x724 ;
  assign n9753 = n9751 ^ x611 ;
  assign n9752 = n9751 ^ x646 ;
  assign n9754 = n9753 ^ n9752 ;
  assign n9757 = ~x1135 & ~n9754 ;
  assign n9758 = n9757 ^ n9752 ;
  assign n9759 = ~x1134 & n9758 ;
  assign n9760 = n9759 ^ n9751 ;
  assign n9764 = n9763 ^ n9760 ;
  assign n9765 = ~x1136 & ~n9764 ;
  assign n9766 = n9765 ^ n9760 ;
  assign n9767 = n9396 & ~n9766 ;
  assign n9768 = ~n9749 & ~n9767 ;
  assign n9798 = x808 ^ x616 ;
  assign n9799 = ~x1136 & n9798 ;
  assign n9800 = n9799 ^ x616 ;
  assign n9802 = n9800 ^ x758 ;
  assign n9801 = n9800 ^ x850 ;
  assign n9803 = n9802 ^ n9801 ;
  assign n9806 = x1136 & n9803 ;
  assign n9807 = n9806 ^ n9801 ;
  assign n9808 = x1134 & n9807 ;
  assign n9809 = n9808 ^ n9800 ;
  assign n9791 = x736 ^ x661 ;
  assign n9792 = n9791 ^ x781 ;
  assign n9795 = x1136 & n9792 ;
  assign n9796 = n9795 ^ x781 ;
  assign n9797 = n9398 & n9796 ;
  assign n9810 = n9809 ^ n9797 ;
  assign n9790 = x736 & x1136 ;
  assign n9811 = n9810 ^ n9790 ;
  assign n9812 = x1135 & n9811 ;
  assign n9813 = n9812 ^ n9809 ;
  assign n9814 = n9395 & n9813 ;
  assign n9769 = x397 ^ x372 ;
  assign n9772 = x592 & n9769 ;
  assign n9773 = n9772 ^ x397 ;
  assign n9774 = n9424 & n9773 ;
  assign n9775 = n9774 ^ x320 ;
  assign n9780 = n9441 & n9775 ;
  assign n9776 = x422 & ~n9436 ;
  assign n9778 = n9776 ^ n9774 ;
  assign n9781 = n9780 ^ n9778 ;
  assign n9815 = n9814 ^ n9781 ;
  assign n9787 = x199 & n7765 ;
  assign n9783 = n9781 ^ x290 ;
  assign n9788 = n9787 ^ n9783 ;
  assign n9789 = ~n9423 & n9788 ;
  assign n9816 = n9815 ^ n9789 ;
  assign n9817 = n3209 & n9816 ;
  assign n9818 = n9817 ^ n9814 ;
  assign n9827 = x866 ^ x749 ;
  assign n9828 = ~x1136 & n9827 ;
  assign n9829 = n9828 ^ x749 ;
  assign n9831 = n9829 ^ x617 ;
  assign n9830 = n9829 ^ x814 ;
  assign n9832 = n9831 ^ n9830 ;
  assign n9835 = x1136 & ~n9832 ;
  assign n9836 = n9835 ^ n9830 ;
  assign n9837 = ~x1134 & ~n9836 ;
  assign n9838 = n9837 ^ n9829 ;
  assign n9820 = x706 ^ x637 ;
  assign n9821 = n9820 ^ x788 ;
  assign n9824 = x1136 & n9821 ;
  assign n9825 = n9824 ^ x788 ;
  assign n9826 = n9398 & n9825 ;
  assign n9839 = n9838 ^ n9826 ;
  assign n9819 = x706 & x1136 ;
  assign n9840 = n9839 ^ n9819 ;
  assign n9841 = x1135 & n9840 ;
  assign n9842 = n9841 ^ n9838 ;
  assign n9843 = n9396 & n9842 ;
  assign n9850 = x411 ^ x387 ;
  assign n9853 = x592 & n9850 ;
  assign n9854 = n9853 ^ x411 ;
  assign n9855 = n9425 & n9854 ;
  assign n9856 = n9855 ^ n9423 ;
  assign n9857 = x452 & n9441 ;
  assign n9858 = n9856 & n9857 ;
  assign n9859 = n9858 ^ x435 ;
  assign n9846 = x199 & n7780 ;
  assign n9847 = n9846 ^ x295 ;
  assign n9848 = n9443 & ~n9847 ;
  assign n9849 = n9848 ^ n3209 ;
  assign n9860 = n9858 ^ n9856 ;
  assign n9861 = n9849 & n9860 ;
  assign n9862 = ~n9436 & n9861 ;
  assign n9863 = n9859 & n9862 ;
  assign n9864 = n9863 ^ n9861 ;
  assign n9865 = n9864 ^ n9849 ;
  assign n9866 = ~n9843 & ~n9865 ;
  assign n9896 = x804 ^ x622 ;
  assign n9897 = ~x1136 & n9896 ;
  assign n9898 = n9897 ^ x622 ;
  assign n9900 = n9898 ^ x743 ;
  assign n9899 = n9898 ^ x859 ;
  assign n9901 = n9900 ^ n9899 ;
  assign n9904 = x1136 & n9901 ;
  assign n9905 = n9904 ^ n9899 ;
  assign n9906 = x1134 & n9905 ;
  assign n9907 = n9906 ^ n9898 ;
  assign n9889 = x735 ^ x639 ;
  assign n9890 = n9889 ^ x783 ;
  assign n9893 = x1136 & n9890 ;
  assign n9894 = n9893 ^ x783 ;
  assign n9895 = n9398 & n9894 ;
  assign n9908 = n9907 ^ n9895 ;
  assign n9888 = x735 & x1136 ;
  assign n9909 = n9908 ^ n9888 ;
  assign n9910 = x1135 & n9909 ;
  assign n9911 = n9910 ^ n9907 ;
  assign n9912 = n9395 & n9911 ;
  assign n9867 = x463 ^ x336 ;
  assign n9870 = x592 & n9867 ;
  assign n9871 = n9870 ^ x463 ;
  assign n9872 = n9424 & n9871 ;
  assign n9873 = n9872 ^ x362 ;
  assign n9878 = n9441 & n9873 ;
  assign n9874 = x437 & ~n9436 ;
  assign n9876 = n9874 ^ n9872 ;
  assign n9879 = n9878 ^ n9876 ;
  assign n9913 = n9912 ^ n9879 ;
  assign n9881 = n9879 ^ x256 ;
  assign n9880 = n9879 ^ x1070 ;
  assign n9882 = n9881 ^ n9880 ;
  assign n9885 = x199 & n9882 ;
  assign n9886 = n9885 ^ n9881 ;
  assign n9887 = ~n9423 & n9886 ;
  assign n9914 = n9913 ^ n9887 ;
  assign n9915 = n3209 & n9914 ;
  assign n9916 = n9915 ^ n9912 ;
  assign n9925 = x803 ^ x623 ;
  assign n9926 = ~x1136 & ~n9925 ;
  assign n9927 = n9926 ^ x623 ;
  assign n9929 = n9927 ^ x748 ;
  assign n9928 = n9927 ^ x876 ;
  assign n9930 = n9929 ^ n9928 ;
  assign n9933 = x1136 & n9930 ;
  assign n9934 = n9933 ^ n9928 ;
  assign n9935 = x1134 & n9934 ;
  assign n9936 = n9935 ^ n9927 ;
  assign n9918 = x730 ^ x710 ;
  assign n9919 = n9918 ^ x789 ;
  assign n9922 = x1136 & n9919 ;
  assign n9923 = n9922 ^ x789 ;
  assign n9924 = n9398 & n9923 ;
  assign n9937 = n9936 ^ n9924 ;
  assign n9917 = x730 & x1136 ;
  assign n9938 = n9937 ^ n9917 ;
  assign n9939 = x1135 & n9938 ;
  assign n9940 = n9939 ^ n9936 ;
  assign n9941 = n9396 & n9940 ;
  assign n9948 = x412 ^ x388 ;
  assign n9951 = x592 & n9948 ;
  assign n9952 = n9951 ^ x412 ;
  assign n9953 = n9425 & n9952 ;
  assign n9954 = n9953 ^ n9423 ;
  assign n9955 = x455 & n9441 ;
  assign n9956 = n9954 & n9955 ;
  assign n9957 = n9956 ^ x436 ;
  assign n9944 = x199 & n7783 ;
  assign n9945 = n9944 ^ x296 ;
  assign n9946 = n9443 & ~n9945 ;
  assign n9947 = n9946 ^ n3209 ;
  assign n9958 = n9956 ^ n9954 ;
  assign n9959 = n9947 & n9958 ;
  assign n9960 = ~n9436 & n9959 ;
  assign n9961 = n9957 & n9960 ;
  assign n9962 = n9961 ^ n9959 ;
  assign n9963 = n9962 ^ n9947 ;
  assign n9964 = ~n9941 & ~n9963 ;
  assign n9994 = x881 ^ x746 ;
  assign n9995 = ~x1136 & n9994 ;
  assign n9996 = n9995 ^ x746 ;
  assign n9998 = n9996 ^ x606 ;
  assign n9997 = n9996 ^ x812 ;
  assign n9999 = n9998 ^ n9997 ;
  assign n10002 = x1136 & ~n9999 ;
  assign n10003 = n10002 ^ n9997 ;
  assign n10004 = ~x1134 & ~n10003 ;
  assign n10005 = n10004 ^ n9996 ;
  assign n9987 = x729 ^ x643 ;
  assign n9988 = n9987 ^ x787 ;
  assign n9991 = x1136 & n9988 ;
  assign n9992 = n9991 ^ x787 ;
  assign n9993 = n9398 & n9992 ;
  assign n10006 = n10005 ^ n9993 ;
  assign n9986 = x729 & x1136 ;
  assign n10007 = n10006 ^ n9986 ;
  assign n10008 = x1135 & n10007 ;
  assign n10009 = n10008 ^ n10005 ;
  assign n10010 = n9395 & n10009 ;
  assign n9965 = x410 ^ x386 ;
  assign n9968 = x592 & n9965 ;
  assign n9969 = n9968 ^ x410 ;
  assign n9970 = n9424 & n9969 ;
  assign n9971 = n9970 ^ x361 ;
  assign n9976 = n9441 & n9971 ;
  assign n9972 = x434 & ~n9436 ;
  assign n9974 = n9972 ^ n9970 ;
  assign n9977 = n9976 ^ n9974 ;
  assign n10011 = n10010 ^ n9977 ;
  assign n9983 = x199 & n7774 ;
  assign n9979 = n9977 ^ x293 ;
  assign n9984 = n9983 ^ n9979 ;
  assign n9985 = ~n9423 & n9984 ;
  assign n10012 = n10011 ^ n9985 ;
  assign n10013 = n3209 & n10012 ;
  assign n10014 = n10013 ^ n10010 ;
  assign n10033 = x366 ^ x335 ;
  assign n10036 = ~x592 & n10033 ;
  assign n10037 = n10036 ^ x366 ;
  assign n10038 = n9424 & n10037 ;
  assign n10039 = n10038 ^ x344 ;
  assign n10044 = n9441 & n10039 ;
  assign n10040 = x416 & ~n9436 ;
  assign n10042 = n10040 ^ n10038 ;
  assign n10045 = n10044 ^ n10042 ;
  assign n10047 = n10045 ^ x259 ;
  assign n10046 = n10045 ^ x1069 ;
  assign n10048 = n10047 ^ n10046 ;
  assign n10051 = x199 & n10048 ;
  assign n10052 = n10051 ^ n10047 ;
  assign n10053 = ~n9423 & n10052 ;
  assign n10054 = n10053 ^ n10045 ;
  assign n10028 = x870 & n9678 ;
  assign n6004 = x742 ^ x704 ;
  assign n10015 = ~x1135 & n6004 ;
  assign n10016 = n10015 ^ x704 ;
  assign n10018 = n10016 ^ x620 ;
  assign n10017 = n10016 ^ x635 ;
  assign n10019 = n10018 ^ n10017 ;
  assign n10022 = ~x1135 & ~n10019 ;
  assign n10023 = n10022 ^ n10017 ;
  assign n10024 = ~x1134 & n10023 ;
  assign n10025 = n10024 ^ n10016 ;
  assign n10029 = n10028 ^ n10025 ;
  assign n10030 = ~x1136 & ~n10029 ;
  assign n10031 = n10030 ^ n10025 ;
  assign n10032 = n9395 & ~n10031 ;
  assign n10055 = n10054 ^ n10032 ;
  assign n10056 = ~n3209 & n10055 ;
  assign n10057 = n10056 ^ n10054 ;
  assign n10071 = x856 & n9678 ;
  assign n6038 = x760 ^ x688 ;
  assign n10058 = ~x1135 & n6038 ;
  assign n10059 = n10058 ^ x688 ;
  assign n10061 = n10059 ^ x613 ;
  assign n10060 = n10059 ^ x632 ;
  assign n10062 = n10061 ^ n10060 ;
  assign n10065 = ~x1135 & ~n10062 ;
  assign n10066 = n10065 ^ n10060 ;
  assign n10067 = ~x1134 & n10066 ;
  assign n10068 = n10067 ^ n10059 ;
  assign n10072 = n10071 ^ n10068 ;
  assign n10073 = ~x1136 & ~n10072 ;
  assign n10074 = n10073 ^ n10068 ;
  assign n10075 = n9396 & ~n10074 ;
  assign n10076 = x1067 ^ x260 ;
  assign n10079 = x199 & n10076 ;
  assign n10080 = n10079 ^ x260 ;
  assign n10081 = n9443 & ~n10080 ;
  assign n10082 = n10081 ^ n3209 ;
  assign n10102 = x346 & n9441 ;
  assign n10103 = n10102 ^ x346 ;
  assign n10083 = x393 & ~x590 ;
  assign n10084 = ~x592 & n10083 ;
  assign n10085 = n10084 ^ x368 ;
  assign n10088 = n10084 ^ x590 ;
  assign n10089 = ~x591 & ~n10088 ;
  assign n10090 = n10085 & n10089 ;
  assign n10091 = n10090 ^ n10085 ;
  assign n10092 = n10091 ^ x368 ;
  assign n10093 = n9435 & ~n10092 ;
  assign n10094 = n10093 ^ n9435 ;
  assign n10095 = n10094 ^ x346 ;
  assign n10104 = n10103 ^ n10095 ;
  assign n10105 = n9423 & ~n10104 ;
  assign n10106 = n10082 & n10105 ;
  assign n10114 = x418 & n10106 ;
  assign n10115 = ~n9436 & n10114 ;
  assign n10116 = n10115 ^ n9436 ;
  assign n10107 = n10106 ^ n10082 ;
  assign n10108 = n10107 ^ n9436 ;
  assign n10117 = n10116 ^ n10108 ;
  assign n10118 = ~n10075 & ~n10117 ;
  assign n10127 = x810 ^ x621 ;
  assign n10128 = ~x1136 & n10127 ;
  assign n10129 = n10128 ^ x621 ;
  assign n10131 = n10129 ^ x739 ;
  assign n10130 = n10129 ^ x874 ;
  assign n10132 = n10131 ^ n10130 ;
  assign n10135 = x1136 & n10132 ;
  assign n10136 = n10135 ^ n10130 ;
  assign n10137 = x1134 & n10136 ;
  assign n10138 = n10137 ^ n10129 ;
  assign n10120 = x690 ^ x665 ;
  assign n10121 = n10120 ^ x791 ;
  assign n10124 = x1136 & n10121 ;
  assign n10125 = n10124 ^ x791 ;
  assign n10126 = n9398 & n10125 ;
  assign n10139 = n10138 ^ n10126 ;
  assign n10119 = x690 & x1136 ;
  assign n10140 = n10139 ^ n10119 ;
  assign n10141 = x1135 & n10140 ;
  assign n10142 = n10141 ^ n10138 ;
  assign n10143 = n9396 & n10142 ;
  assign n10144 = x413 ^ x389 ;
  assign n10147 = x592 & n10144 ;
  assign n10148 = n10147 ^ x413 ;
  assign n10149 = n9425 & n10148 ;
  assign n10150 = n10149 ^ n9423 ;
  assign n10151 = x450 & n9441 ;
  assign n10152 = n10150 & n10151 ;
  assign n10153 = n10152 ^ x438 ;
  assign n10154 = n10152 ^ n10150 ;
  assign n10155 = x1036 ^ x255 ;
  assign n10158 = x199 & n10155 ;
  assign n10159 = n10158 ^ x255 ;
  assign n10160 = n9443 & ~n10159 ;
  assign n10161 = n10160 ^ n3209 ;
  assign n10162 = n10154 & n10161 ;
  assign n10163 = ~n9436 & n10162 ;
  assign n10164 = n10153 & n10163 ;
  assign n10165 = n10164 ^ n10162 ;
  assign n10166 = n10165 ^ n10161 ;
  assign n10167 = ~n10143 & ~n10166 ;
  assign n10168 = x1100 ^ x680 ;
  assign n10171 = n9163 & n10168 ;
  assign n10172 = n10171 ^ x680 ;
  assign n10173 = ~x962 & n10172 ;
  assign n10174 = x1103 ^ x681 ;
  assign n10177 = n9163 & n10174 ;
  assign n10178 = n10177 ^ x681 ;
  assign n10179 = ~x962 & n10178 ;
  assign n10180 = x392 ^ x367 ;
  assign n10183 = x592 & n10180 ;
  assign n10184 = n10183 ^ x392 ;
  assign n10185 = n9425 & n10184 ;
  assign n10186 = n10185 ^ n9423 ;
  assign n10187 = x417 & ~n9436 ;
  assign n10188 = n10186 & n10187 ;
  assign n10189 = n10188 ^ x345 ;
  assign n10190 = n10188 ^ n10186 ;
  assign n10191 = x1039 ^ x251 ;
  assign n10194 = x199 & n10191 ;
  assign n10195 = n10194 ^ x251 ;
  assign n10196 = n9443 & ~n10195 ;
  assign n10197 = n10196 ^ n3209 ;
  assign n10198 = n10190 & n10197 ;
  assign n10199 = n9441 & n10198 ;
  assign n10200 = n10189 & n10199 ;
  assign n10201 = n10200 ^ n10198 ;
  assign n10202 = n10201 ^ n10197 ;
  assign n10216 = x848 & n9678 ;
  assign n6016 = x757 ^ x686 ;
  assign n10203 = ~x1135 & n6016 ;
  assign n10204 = n10203 ^ x686 ;
  assign n10206 = n10204 ^ x610 ;
  assign n10205 = n10204 ^ x631 ;
  assign n10207 = n10206 ^ n10205 ;
  assign n10210 = ~x1135 & ~n10207 ;
  assign n10211 = n10210 ^ n10205 ;
  assign n10212 = ~x1134 & n10211 ;
  assign n10213 = n10212 ^ n10204 ;
  assign n10217 = n10216 ^ n10213 ;
  assign n10218 = ~x1136 & ~n10217 ;
  assign n10219 = n10218 ^ n10213 ;
  assign n10220 = n9396 & ~n10219 ;
  assign n10221 = ~n10202 & ~n10220 ;
  assign n10222 = x1130 ^ x684 ;
  assign n10225 = n9162 & ~n10222 ;
  assign n10226 = n10225 ^ x684 ;
  assign n10227 = ~x962 & ~n10226 ;
  assign n10234 = x744 ^ x728 ;
  assign n10235 = ~x1135 & n10234 ;
  assign n10236 = n10235 ^ x728 ;
  assign n10238 = n10236 ^ x652 ;
  assign n10237 = n10236 ^ x657 ;
  assign n10239 = n10238 ^ n10237 ;
  assign n10242 = ~x1135 & ~n10239 ;
  assign n10243 = n10242 ^ n10237 ;
  assign n10244 = ~x1134 & n10243 ;
  assign n10245 = n10244 ^ n10236 ;
  assign n10228 = x860 ^ x813 ;
  assign n10231 = ~x1134 & n10228 ;
  assign n10232 = n10231 ^ x860 ;
  assign n10233 = ~x1135 & n10232 ;
  assign n10246 = n10245 ^ n10233 ;
  assign n10247 = ~x1136 & ~n10246 ;
  assign n10248 = n10247 ^ n10245 ;
  assign n10249 = n9396 & ~n10248 ;
  assign n10250 = x406 ^ x382 ;
  assign n10253 = x592 & n10250 ;
  assign n10254 = n10253 ^ x406 ;
  assign n10255 = n9425 & n10254 ;
  assign n10256 = n10255 ^ n9423 ;
  assign n10257 = x430 & ~n9436 ;
  assign n10258 = n10256 & n10257 ;
  assign n10259 = n10258 ^ x357 ;
  assign n10260 = n10258 ^ n10256 ;
  assign n10261 = n7480 ^ x1076 ;
  assign n10264 = ~x199 & n10261 ;
  assign n10265 = n10264 ^ x1076 ;
  assign n10266 = n9443 & ~n10265 ;
  assign n10267 = n10266 ^ n3209 ;
  assign n10268 = n10260 & n10267 ;
  assign n10269 = n9441 & n10268 ;
  assign n10270 = n10259 & n10269 ;
  assign n10271 = n10270 ^ n10268 ;
  assign n10272 = n10271 ^ n10267 ;
  assign n10273 = ~n10249 & ~n10272 ;
  assign n10274 = x1113 ^ x686 ;
  assign n10277 = n9162 & ~n10274 ;
  assign n10278 = n10277 ^ x686 ;
  assign n10279 = ~x962 & ~n10278 ;
  assign n10280 = x1127 ^ x687 ;
  assign n10283 = n9162 & n10280 ;
  assign n10284 = n10283 ^ x687 ;
  assign n10285 = ~x962 & n10284 ;
  assign n10286 = x1115 ^ x688 ;
  assign n10289 = n9162 & ~n10286 ;
  assign n10290 = n10289 ^ x688 ;
  assign n10291 = ~x962 & ~n10290 ;
  assign n6112 = x752 ^ x703 ;
  assign n10319 = ~x1135 & ~n6112 ;
  assign n10320 = n10319 ^ x703 ;
  assign n10322 = n10320 ^ x655 ;
  assign n10321 = n10320 ^ x658 ;
  assign n10323 = n10322 ^ n10321 ;
  assign n10326 = x1135 & ~n10323 ;
  assign n10327 = n10326 ^ n10321 ;
  assign n10328 = ~x1134 & n10327 ;
  assign n10329 = n10328 ^ n10320 ;
  assign n10313 = x843 ^ x798 ;
  assign n10316 = ~x1134 & n10313 ;
  assign n10317 = n10316 ^ x843 ;
  assign n10318 = ~x1135 & n10317 ;
  assign n10330 = n10329 ^ n10318 ;
  assign n10331 = ~x1136 & n10330 ;
  assign n10332 = n10331 ^ n10329 ;
  assign n10333 = n9395 & n10332 ;
  assign n10292 = x401 ^ x376 ;
  assign n10295 = x592 & n10292 ;
  assign n10296 = n10295 ^ x401 ;
  assign n10297 = n9424 & n10296 ;
  assign n10298 = n10297 ^ x351 ;
  assign n10303 = n9441 & n10298 ;
  assign n10299 = x426 & ~n9436 ;
  assign n10301 = n10299 ^ n10297 ;
  assign n10304 = n10303 ^ n10301 ;
  assign n10334 = n10333 ^ n10304 ;
  assign n10306 = n10304 ^ x1079 ;
  assign n10305 = n10304 ^ n7450 ;
  assign n10307 = n10306 ^ n10305 ;
  assign n10310 = ~x199 & n10307 ;
  assign n10311 = n10310 ^ n10306 ;
  assign n10312 = ~n9423 & n10311 ;
  assign n10335 = n10334 ^ n10312 ;
  assign n10336 = n3209 & n10335 ;
  assign n10337 = n10336 ^ n10333 ;
  assign n10338 = x1108 ^ x690 ;
  assign n10341 = n9162 & n10338 ;
  assign n10342 = n10341 ^ x690 ;
  assign n10343 = ~x962 & n10342 ;
  assign n10344 = x1107 ^ x691 ;
  assign n10347 = n9162 & n10344 ;
  assign n10348 = n10347 ^ x691 ;
  assign n10349 = ~x962 & n10348 ;
  assign n5912 = x770 ^ x726 ;
  assign n10356 = ~x1135 & ~n5912 ;
  assign n10357 = n10356 ^ x726 ;
  assign n10359 = n10357 ^ x649 ;
  assign n10358 = n10357 ^ x656 ;
  assign n10360 = n10359 ^ n10358 ;
  assign n10363 = x1135 & ~n10360 ;
  assign n10364 = n10363 ^ n10358 ;
  assign n10365 = ~x1134 & n10364 ;
  assign n10366 = n10365 ^ n10357 ;
  assign n10350 = x844 ^ x801 ;
  assign n10353 = ~x1134 & n10350 ;
  assign n10354 = n10353 ^ x844 ;
  assign n10355 = ~x1135 & n10354 ;
  assign n10367 = n10366 ^ n10355 ;
  assign n10368 = ~x1136 & n10367 ;
  assign n10369 = n10368 ^ n10366 ;
  assign n10370 = n9396 & n10369 ;
  assign n10371 = x402 ^ x317 ;
  assign n10374 = x592 & n10371 ;
  assign n10375 = n10374 ^ x402 ;
  assign n10376 = n9425 & n10375 ;
  assign n10377 = n10376 ^ n9423 ;
  assign n10378 = x427 & ~n9436 ;
  assign n10379 = n10377 & n10378 ;
  assign n10380 = n10379 ^ x352 ;
  assign n10381 = n10379 ^ n10377 ;
  assign n10382 = n7462 ^ x1078 ;
  assign n10385 = ~x199 & n10382 ;
  assign n10386 = n10385 ^ x1078 ;
  assign n10387 = n9443 & ~n10386 ;
  assign n10388 = n10387 ^ n3209 ;
  assign n10389 = n10381 & n10388 ;
  assign n10390 = n9441 & n10389 ;
  assign n10391 = n10380 & n10390 ;
  assign n10392 = n10391 ^ n10389 ;
  assign n10393 = n10392 ^ n10388 ;
  assign n10394 = ~n10370 & ~n10393 ;
  assign n10395 = x1129 ^ x693 ;
  assign n10398 = n9163 & ~n10395 ;
  assign n10399 = n10398 ^ x693 ;
  assign n10400 = ~x962 & ~n10399 ;
  assign n10401 = x1128 ^ x694 ;
  assign n10404 = n9162 & ~n10401 ;
  assign n10405 = n10404 ^ x694 ;
  assign n10406 = ~x962 & ~n10405 ;
  assign n10407 = x1111 ^ x695 ;
  assign n10410 = n9163 & ~n10407 ;
  assign n10411 = n10410 ^ x695 ;
  assign n10412 = ~x962 & ~n10411 ;
  assign n10413 = x1100 ^ x696 ;
  assign n10416 = n9162 & n10413 ;
  assign n10417 = n10416 ^ x696 ;
  assign n10418 = ~x962 & n10417 ;
  assign n10419 = x1129 ^ x697 ;
  assign n10422 = n9162 & ~n10419 ;
  assign n10423 = n10422 ^ x697 ;
  assign n10424 = ~x962 & ~n10423 ;
  assign n10425 = x1116 ^ x698 ;
  assign n10428 = n9162 & ~n10425 ;
  assign n10429 = n10428 ^ x698 ;
  assign n10430 = ~x962 & ~n10429 ;
  assign n10431 = x1103 ^ x699 ;
  assign n10434 = n9162 & n10431 ;
  assign n10435 = n10434 ^ x699 ;
  assign n10436 = ~x962 & n10435 ;
  assign n10437 = x1110 ^ x700 ;
  assign n10440 = n9162 & n10437 ;
  assign n10441 = n10440 ^ x700 ;
  assign n10442 = ~x962 & n10441 ;
  assign n10443 = x1123 ^ x701 ;
  assign n10446 = n9162 & ~n10443 ;
  assign n10447 = n10446 ^ x701 ;
  assign n10448 = ~x962 & ~n10447 ;
  assign n10449 = x1117 ^ x702 ;
  assign n10452 = n9162 & ~n10449 ;
  assign n10453 = n10452 ^ x702 ;
  assign n10454 = ~x962 & ~n10453 ;
  assign n10455 = x1124 ^ x703 ;
  assign n10458 = n9162 & n10455 ;
  assign n10459 = n10458 ^ x703 ;
  assign n10460 = ~x962 & n10459 ;
  assign n10461 = x1112 ^ x704 ;
  assign n10464 = n9162 & ~n10461 ;
  assign n10465 = n10464 ^ x704 ;
  assign n10466 = ~x962 & ~n10465 ;
  assign n10467 = x1125 ^ x705 ;
  assign n10470 = n9162 & n10467 ;
  assign n10471 = n10470 ^ x705 ;
  assign n10472 = ~x962 & n10471 ;
  assign n10473 = x1105 ^ x706 ;
  assign n10476 = n9162 & n10473 ;
  assign n10477 = n10476 ^ x706 ;
  assign n10478 = ~x962 & n10477 ;
  assign n10479 = x395 ^ x370 ;
  assign n10482 = x592 & n10479 ;
  assign n10483 = n10482 ^ x395 ;
  assign n10484 = n9425 & n10483 ;
  assign n10485 = n10484 ^ n9423 ;
  assign n10486 = x420 & ~n9436 ;
  assign n10487 = n10485 & n10486 ;
  assign n10488 = n10487 ^ x347 ;
  assign n10494 = x200 & n7833 ;
  assign n10490 = x1055 ^ x304 ;
  assign n10495 = n10494 ^ n10490 ;
  assign n10496 = ~x199 & n10495 ;
  assign n10497 = n10496 ^ x1055 ;
  assign n10498 = ~n9423 & ~n10497 ;
  assign n10499 = n3209 & ~n10498 ;
  assign n10500 = n10487 ^ n10485 ;
  assign n10501 = n10499 & n10500 ;
  assign n10502 = n9441 & n10501 ;
  assign n10503 = n10488 & n10502 ;
  assign n10504 = n10503 ^ n10501 ;
  assign n10505 = n10504 ^ n10499 ;
  assign n10519 = x847 & n9678 ;
  assign n6051 = x753 ^ x702 ;
  assign n10506 = ~x1135 & n6051 ;
  assign n10507 = n10506 ^ x702 ;
  assign n10509 = n10507 ^ x618 ;
  assign n10508 = n10507 ^ x627 ;
  assign n10510 = n10509 ^ n10508 ;
  assign n10513 = ~x1135 & n10510 ;
  assign n10514 = n10513 ^ n10508 ;
  assign n10515 = ~x1134 & ~n10514 ;
  assign n10516 = n10515 ^ n10507 ;
  assign n10520 = n10519 ^ n10516 ;
  assign n10521 = ~x1136 & ~n10520 ;
  assign n10522 = n10521 ^ n10516 ;
  assign n10523 = n9396 & ~n10522 ;
  assign n10524 = ~n10505 & ~n10523 ;
  assign n10551 = x442 ^ x328 ;
  assign n10554 = ~x592 & n10551 ;
  assign n10555 = n10554 ^ x442 ;
  assign n10556 = n9424 & n10555 ;
  assign n10557 = n10556 ^ x321 ;
  assign n10562 = n9441 & n10557 ;
  assign n10558 = x459 & ~n9436 ;
  assign n10560 = n10558 ^ n10556 ;
  assign n10563 = n10562 ^ n10560 ;
  assign n10564 = n10563 ^ x1058 ;
  assign n10548 = x200 & n7836 ;
  assign n10544 = x1058 ^ x305 ;
  assign n10549 = n10548 ^ n10544 ;
  assign n10550 = ~x199 & n10549 ;
  assign n10565 = n10564 ^ n10550 ;
  assign n10566 = ~n9423 & n10565 ;
  assign n10567 = n10566 ^ n10563 ;
  assign n10538 = x857 & n9678 ;
  assign n6061 = x754 ^ x709 ;
  assign n10525 = ~x1135 & n6061 ;
  assign n10526 = n10525 ^ x709 ;
  assign n10528 = n10526 ^ x609 ;
  assign n10527 = n10526 ^ x660 ;
  assign n10529 = n10528 ^ n10527 ;
  assign n10532 = ~x1135 & n10529 ;
  assign n10533 = n10532 ^ n10527 ;
  assign n10534 = ~x1134 & ~n10533 ;
  assign n10535 = n10534 ^ n10526 ;
  assign n10539 = n10538 ^ n10535 ;
  assign n10540 = ~x1136 & ~n10539 ;
  assign n10541 = n10540 ^ n10535 ;
  assign n10542 = n9395 & ~n10541 ;
  assign n10568 = n10567 ^ n10542 ;
  assign n10569 = ~n3209 & n10568 ;
  assign n10570 = n10569 ^ n10567 ;
  assign n10571 = x1118 ^ x709 ;
  assign n10574 = n9162 & ~n10571 ;
  assign n10575 = n10574 ^ x709 ;
  assign n10576 = ~x962 & ~n10575 ;
  assign n10577 = x1106 ^ x710 ;
  assign n10580 = n9163 & n10577 ;
  assign n10581 = n10580 ^ x710 ;
  assign n10582 = ~x962 & n10581 ;
  assign n10583 = x398 ^ x373 ;
  assign n10586 = x592 & n10583 ;
  assign n10587 = n10586 ^ x398 ;
  assign n10588 = n9425 & n10587 ;
  assign n10589 = n10588 ^ n9423 ;
  assign n10590 = x423 & ~n9436 ;
  assign n10591 = n10589 & n10590 ;
  assign n10592 = n10591 ^ x348 ;
  assign n10598 = x200 & n7839 ;
  assign n10594 = x1087 ^ x306 ;
  assign n10599 = n10598 ^ n10594 ;
  assign n10600 = ~x199 & n10599 ;
  assign n10601 = n10600 ^ x1087 ;
  assign n10602 = ~n9423 & ~n10601 ;
  assign n10603 = n3209 & ~n10602 ;
  assign n10604 = n10591 ^ n10589 ;
  assign n10605 = n10603 & n10604 ;
  assign n10606 = n9441 & n10605 ;
  assign n10607 = n10592 & n10606 ;
  assign n10608 = n10607 ^ n10605 ;
  assign n10609 = n10608 ^ n10603 ;
  assign n10623 = x858 & n9678 ;
  assign n5947 = x755 ^ x725 ;
  assign n10610 = ~x1135 & n5947 ;
  assign n10611 = n10610 ^ x725 ;
  assign n10613 = n10611 ^ x630 ;
  assign n10612 = n10611 ^ x647 ;
  assign n10614 = n10613 ^ n10612 ;
  assign n10617 = ~x1135 & n10614 ;
  assign n10618 = n10617 ^ n10612 ;
  assign n10619 = ~x1134 & ~n10618 ;
  assign n10620 = n10619 ^ n10611 ;
  assign n10624 = n10623 ^ n10620 ;
  assign n10625 = ~x1136 & ~n10624 ;
  assign n10626 = n10625 ^ n10620 ;
  assign n10627 = n9396 & ~n10626 ;
  assign n10628 = ~n10609 & ~n10627 ;
  assign n10629 = x400 ^ x374 ;
  assign n10632 = x592 & n10629 ;
  assign n10633 = n10632 ^ x400 ;
  assign n10634 = n9425 & n10633 ;
  assign n10635 = n10634 ^ n9423 ;
  assign n10636 = x425 & ~n9436 ;
  assign n10637 = n10635 & n10636 ;
  assign n10638 = n10637 ^ x350 ;
  assign n10644 = x200 & n7789 ;
  assign n10640 = x1035 ^ x298 ;
  assign n10645 = n10644 ^ n10640 ;
  assign n10646 = ~x199 & n10645 ;
  assign n10647 = n10646 ^ x1035 ;
  assign n10648 = ~n9423 & ~n10647 ;
  assign n10649 = n3209 & ~n10648 ;
  assign n10650 = n10637 ^ n10635 ;
  assign n10651 = n10649 & n10650 ;
  assign n10652 = n9441 & n10651 ;
  assign n10653 = n10638 & n10652 ;
  assign n10654 = n10653 ^ n10651 ;
  assign n10655 = n10654 ^ n10649 ;
  assign n10669 = x842 & n9678 ;
  assign n5959 = x751 ^ x701 ;
  assign n10656 = ~x1135 & n5959 ;
  assign n10657 = n10656 ^ x701 ;
  assign n10659 = n10657 ^ x644 ;
  assign n10658 = n10657 ^ x715 ;
  assign n10660 = n10659 ^ n10658 ;
  assign n10663 = ~x1135 & n10660 ;
  assign n10664 = n10663 ^ n10658 ;
  assign n10665 = ~x1134 & ~n10664 ;
  assign n10666 = n10665 ^ n10657 ;
  assign n10670 = n10669 ^ n10666 ;
  assign n10671 = ~x1136 & ~n10670 ;
  assign n10672 = n10671 ^ n10666 ;
  assign n10673 = n9396 & ~n10672 ;
  assign n10674 = ~n10655 & ~n10673 ;
  assign n10675 = x396 ^ x371 ;
  assign n10678 = x592 & n10675 ;
  assign n10679 = n10678 ^ x396 ;
  assign n10680 = n9425 & n10679 ;
  assign n10681 = n10680 ^ n9423 ;
  assign n10682 = x421 & ~n9436 ;
  assign n10683 = n10681 & n10682 ;
  assign n10684 = n10683 ^ x322 ;
  assign n10690 = x200 & n7848 ;
  assign n10686 = x1051 ^ x309 ;
  assign n10691 = n10690 ^ n10686 ;
  assign n10692 = ~x199 & n10691 ;
  assign n10693 = n10692 ^ x1051 ;
  assign n10694 = ~n9423 & ~n10693 ;
  assign n10695 = n3209 & ~n10694 ;
  assign n10696 = n10683 ^ n10681 ;
  assign n10697 = n10695 & n10696 ;
  assign n10698 = n9441 & n10697 ;
  assign n10699 = n10684 & n10698 ;
  assign n10700 = n10699 ^ n10697 ;
  assign n10701 = n10700 ^ n10695 ;
  assign n10715 = x854 & n9678 ;
  assign n6072 = x756 ^ x734 ;
  assign n10702 = ~x1135 & n6072 ;
  assign n10703 = n10702 ^ x734 ;
  assign n10705 = n10703 ^ x628 ;
  assign n10704 = n10703 ^ x629 ;
  assign n10706 = n10705 ^ n10704 ;
  assign n10709 = x1135 & n10706 ;
  assign n10710 = n10709 ^ n10704 ;
  assign n10711 = ~x1134 & ~n10710 ;
  assign n10712 = n10711 ^ n10703 ;
  assign n10716 = n10715 ^ n10712 ;
  assign n10717 = ~x1136 & ~n10716 ;
  assign n10718 = n10717 ^ n10712 ;
  assign n10719 = n9396 & ~n10718 ;
  assign n10720 = ~n10701 & ~n10719 ;
  assign n10748 = x762 ^ x697 ;
  assign n10749 = ~x1135 & n10748 ;
  assign n10750 = n10749 ^ x697 ;
  assign n10752 = n10750 ^ x653 ;
  assign n10751 = n10750 ^ x693 ;
  assign n10753 = n10752 ^ n10751 ;
  assign n10756 = ~x1135 & ~n10753 ;
  assign n10757 = n10756 ^ n10751 ;
  assign n10758 = ~x1134 & n10757 ;
  assign n10759 = n10758 ^ n10750 ;
  assign n10742 = x867 ^ x816 ;
  assign n10745 = ~x1134 & n10742 ;
  assign n10746 = n10745 ^ x867 ;
  assign n10747 = ~x1135 & n10746 ;
  assign n10760 = n10759 ^ n10747 ;
  assign n10761 = ~x1136 & ~n10760 ;
  assign n10762 = n10761 ^ n10759 ;
  assign n10763 = n9395 & ~n10762 ;
  assign n10721 = x439 ^ x326 ;
  assign n10724 = ~x592 & n10721 ;
  assign n10725 = n10724 ^ x439 ;
  assign n10726 = n9424 & n10725 ;
  assign n10727 = n10726 ^ x449 ;
  assign n10732 = ~n9436 & n10727 ;
  assign n10728 = x461 & n9441 ;
  assign n10730 = n10728 ^ n10726 ;
  assign n10733 = n10732 ^ n10730 ;
  assign n10764 = n10763 ^ n10733 ;
  assign n10735 = n10733 ^ x1057 ;
  assign n10734 = n10733 ^ n7414 ;
  assign n10736 = n10735 ^ n10734 ;
  assign n10739 = ~x199 & n10736 ;
  assign n10740 = n10739 ^ n10735 ;
  assign n10741 = ~n9423 & n10740 ;
  assign n10765 = n10764 ^ n10741 ;
  assign n10766 = n3209 & n10765 ;
  assign n10767 = n10766 ^ n10763 ;
  assign n10768 = x1123 ^ x715 ;
  assign n10771 = n9163 & n10768 ;
  assign n10772 = n10771 ^ x715 ;
  assign n10773 = ~x962 & n10772 ;
  assign n10787 = x845 & n9678 ;
  assign n5803 = x761 ^ x738 ;
  assign n10774 = ~x1135 & n5803 ;
  assign n10775 = n10774 ^ x738 ;
  assign n10777 = n10775 ^ x626 ;
  assign n10776 = n10775 ^ x641 ;
  assign n10778 = n10777 ^ n10776 ;
  assign n10781 = ~x1135 & n10778 ;
  assign n10782 = n10781 ^ n10776 ;
  assign n10783 = ~x1134 & ~n10782 ;
  assign n10784 = n10783 ^ n10775 ;
  assign n10788 = n10787 ^ n10784 ;
  assign n10789 = ~x1136 & ~n10788 ;
  assign n10790 = n10789 ^ n10784 ;
  assign n10791 = n9396 & ~n10790 ;
  assign n10797 = x200 & n7842 ;
  assign n10793 = x1043 ^ x307 ;
  assign n10798 = n10797 ^ n10793 ;
  assign n10799 = ~x199 & n10798 ;
  assign n10800 = n10799 ^ x1043 ;
  assign n10801 = ~n9423 & ~n10800 ;
  assign n10802 = n3209 & ~n10801 ;
  assign n10803 = x440 ^ x329 ;
  assign n10806 = ~x592 & n10803 ;
  assign n10807 = n10806 ^ x440 ;
  assign n10808 = n9425 & n10807 ;
  assign n10809 = n10808 ^ n9423 ;
  assign n10810 = n10802 & n10809 ;
  assign n10811 = x349 & n9441 ;
  assign n10812 = n10810 & n10811 ;
  assign n10813 = n10812 ^ n10810 ;
  assign n10821 = x454 & n10813 ;
  assign n10822 = ~n9436 & n10821 ;
  assign n10823 = n10822 ^ n9436 ;
  assign n10814 = n10813 ^ n10802 ;
  assign n10815 = n10814 ^ n9436 ;
  assign n10824 = n10823 ^ n10815 ;
  assign n10825 = ~n10791 & ~n10824 ;
  assign n6144 = x768 ^ x705 ;
  assign n10853 = ~x1135 & ~n6144 ;
  assign n10854 = n10853 ^ x705 ;
  assign n10856 = n10854 ^ x645 ;
  assign n10855 = n10854 ^ x669 ;
  assign n10857 = n10856 ^ n10855 ;
  assign n10860 = ~x1135 & ~n10857 ;
  assign n10861 = n10860 ^ n10855 ;
  assign n10862 = ~x1134 & ~n10861 ;
  assign n10863 = n10862 ^ n10854 ;
  assign n10847 = x839 ^ x800 ;
  assign n10850 = ~x1134 & n10847 ;
  assign n10851 = n10850 ^ x839 ;
  assign n10852 = ~x1135 & n10851 ;
  assign n10864 = n10863 ^ n10852 ;
  assign n10865 = ~x1136 & n10864 ;
  assign n10866 = n10865 ^ n10863 ;
  assign n10867 = n9395 & n10866 ;
  assign n10826 = x377 ^ x318 ;
  assign n10829 = ~x592 & n10826 ;
  assign n10830 = n10829 ^ x377 ;
  assign n10831 = n9424 & n10830 ;
  assign n10832 = n10831 ^ x448 ;
  assign n10837 = ~n9436 & n10832 ;
  assign n10833 = x462 & n9441 ;
  assign n10835 = n10833 ^ n10831 ;
  assign n10838 = n10837 ^ n10835 ;
  assign n10868 = n10867 ^ n10838 ;
  assign n10840 = n10838 ^ x1074 ;
  assign n10839 = n10838 ^ n7456 ;
  assign n10841 = n10840 ^ n10839 ;
  assign n10844 = ~x199 & n10841 ;
  assign n10845 = n10844 ^ n10840 ;
  assign n10846 = ~n9423 & n10845 ;
  assign n10869 = n10868 ^ n10846 ;
  assign n10870 = n3209 & n10869 ;
  assign n10871 = n10870 ^ n10867 ;
  assign n10873 = x419 & ~n9436 ;
  assign n10872 = x315 & n9441 ;
  assign n10874 = n10873 ^ n10872 ;
  assign n10875 = x394 ^ x369 ;
  assign n10878 = x592 & n10875 ;
  assign n10879 = n10878 ^ x394 ;
  assign n10880 = n9425 & n10879 ;
  assign n10881 = n10880 ^ n9423 ;
  assign n10882 = ~n10874 & n10881 ;
  assign n10888 = x200 & n7830 ;
  assign n10884 = x1080 ^ x303 ;
  assign n10889 = n10888 ^ n10884 ;
  assign n10890 = ~x199 & n10889 ;
  assign n10891 = n10890 ^ x1080 ;
  assign n10892 = ~n9423 & ~n10891 ;
  assign n10893 = n3209 & ~n10892 ;
  assign n10894 = ~n10882 & n10893 ;
  assign n10908 = x853 & n9678 ;
  assign n5892 = x767 ^ x698 ;
  assign n10895 = ~x1135 & n5892 ;
  assign n10896 = n10895 ^ x698 ;
  assign n10898 = n10896 ^ x608 ;
  assign n10897 = n10896 ^ x625 ;
  assign n10899 = n10898 ^ n10897 ;
  assign n10902 = ~x1135 & n10899 ;
  assign n10903 = n10902 ^ n10897 ;
  assign n10904 = ~x1134 & ~n10903 ;
  assign n10905 = n10904 ^ n10896 ;
  assign n10909 = n10908 ^ n10905 ;
  assign n10910 = ~x1136 & ~n10909 ;
  assign n10911 = n10910 ^ n10905 ;
  assign n10912 = n9396 & ~n10911 ;
  assign n10913 = ~n10894 & ~n10912 ;
  assign n5870 = x774 ^ x687 ;
  assign n10941 = ~x1135 & ~n5870 ;
  assign n10942 = n10941 ^ x687 ;
  assign n10944 = n10942 ^ x636 ;
  assign n10943 = n10942 ^ x650 ;
  assign n10945 = n10944 ^ n10943 ;
  assign n10948 = ~x1135 & ~n10945 ;
  assign n10949 = n10948 ^ n10943 ;
  assign n10950 = ~x1134 & ~n10949 ;
  assign n10951 = n10950 ^ n10942 ;
  assign n10935 = x868 ^ x807 ;
  assign n10938 = ~x1134 & n10935 ;
  assign n10939 = n10938 ^ x868 ;
  assign n10940 = ~x1135 & n10939 ;
  assign n10952 = n10951 ^ n10940 ;
  assign n10953 = ~x1136 & n10952 ;
  assign n10954 = n10953 ^ n10951 ;
  assign n10955 = n9395 & n10954 ;
  assign n10914 = x378 ^ x325 ;
  assign n10917 = ~x592 & n10914 ;
  assign n10918 = n10917 ^ x378 ;
  assign n10919 = n9424 & n10918 ;
  assign n10920 = n10919 ^ x353 ;
  assign n10925 = n9441 & n10920 ;
  assign n10921 = x451 & ~n9436 ;
  assign n10923 = n10921 ^ n10919 ;
  assign n10926 = n10925 ^ n10923 ;
  assign n10956 = n10955 ^ n10926 ;
  assign n10928 = n10926 ^ x1063 ;
  assign n10927 = n10926 ^ n7468 ;
  assign n10929 = n10928 ^ n10927 ;
  assign n10932 = ~x199 & n10929 ;
  assign n10933 = n10932 ^ n10928 ;
  assign n10934 = ~n9423 & n10933 ;
  assign n10957 = n10956 ^ n10934 ;
  assign n10958 = n3209 & n10957 ;
  assign n10959 = n10958 ^ n10955 ;
  assign n10987 = x750 ^ x684 ;
  assign n10988 = ~x1135 & n10987 ;
  assign n10989 = n10988 ^ x684 ;
  assign n10991 = n10989 ^ x651 ;
  assign n10990 = n10989 ^ x654 ;
  assign n10992 = n10991 ^ n10990 ;
  assign n10995 = ~x1135 & ~n10992 ;
  assign n10996 = n10995 ^ n10990 ;
  assign n10997 = ~x1134 & n10996 ;
  assign n10998 = n10997 ^ n10989 ;
  assign n10981 = x880 ^ x794 ;
  assign n10984 = ~x1134 & n10981 ;
  assign n10985 = n10984 ^ x880 ;
  assign n10986 = ~x1135 & n10985 ;
  assign n10999 = n10998 ^ n10986 ;
  assign n11000 = ~x1136 & ~n10999 ;
  assign n11001 = n11000 ^ n10998 ;
  assign n11002 = n9395 & ~n11001 ;
  assign n10960 = x405 ^ x381 ;
  assign n10963 = x592 & n10960 ;
  assign n10964 = n10963 ^ x405 ;
  assign n10965 = n9424 & n10964 ;
  assign n10966 = n10965 ^ x356 ;
  assign n10971 = n9441 & n10966 ;
  assign n10967 = x445 & ~n9436 ;
  assign n10969 = n10967 ^ n10965 ;
  assign n10972 = n10971 ^ n10969 ;
  assign n11003 = n11002 ^ n10972 ;
  assign n10974 = n10972 ^ x1081 ;
  assign n10973 = n10972 ^ n7486 ;
  assign n10975 = n10974 ^ n10973 ;
  assign n10978 = ~x199 & n10975 ;
  assign n10979 = n10978 ^ n10974 ;
  assign n10980 = ~n9423 & n10979 ;
  assign n11004 = n11003 ^ n10980 ;
  assign n11005 = n3209 & n11004 ;
  assign n11006 = n11005 ^ n11002 ;
  assign n11007 = x807 ^ x747 ;
  assign n11008 = x798 ^ x765 ;
  assign n11009 = x800 ^ x771 ;
  assign n11010 = ~n11008 & ~n11009 ;
  assign n11011 = x816 ^ x775 ;
  assign n11012 = n11010 & ~n11011 ;
  assign n11013 = ~n11007 & n11012 ;
  assign n11014 = x813 ^ x721 ;
  assign n11015 = x794 ^ x769 ;
  assign n11016 = x801 ^ x773 ;
  assign n11017 = ~n11015 & ~n11016 ;
  assign n11018 = x795 ^ x731 ;
  assign n11019 = n11017 & ~n11018 ;
  assign n11020 = ~n11014 & n11019 ;
  assign n11021 = n11013 & n11020 ;
  assign n11022 = x747 & x773 ;
  assign n11023 = x731 & ~x945 ;
  assign n11024 = n11022 & n11023 ;
  assign n11025 = x775 & x988 ;
  assign n11026 = n11024 & n11025 ;
  assign n11031 = x769 & n11026 ;
  assign n11032 = n11031 ^ x721 ;
  assign n11033 = ~n11021 & n11032 ;
  assign n11040 = x776 ^ x694 ;
  assign n11041 = ~x1135 & n11040 ;
  assign n11042 = n11041 ^ x694 ;
  assign n11044 = n11042 ^ x640 ;
  assign n11043 = n11042 ^ x732 ;
  assign n11045 = n11044 ^ n11043 ;
  assign n11048 = ~x1135 & ~n11045 ;
  assign n11049 = n11048 ^ n11043 ;
  assign n11050 = ~x1134 & n11049 ;
  assign n11051 = n11050 ^ n11042 ;
  assign n11034 = x851 ^ x795 ;
  assign n11037 = ~x1134 & n11034 ;
  assign n11038 = n11037 ^ x851 ;
  assign n11039 = ~x1135 & n11038 ;
  assign n11052 = n11051 ^ n11039 ;
  assign n11053 = ~x1136 & ~n11052 ;
  assign n11054 = n11053 ^ n11051 ;
  assign n11055 = n9396 & ~n11054 ;
  assign n11056 = x403 ^ x379 ;
  assign n11059 = x592 & n11056 ;
  assign n11060 = n11059 ^ x403 ;
  assign n11061 = n9425 & n11060 ;
  assign n11062 = n11061 ^ n9423 ;
  assign n11063 = x428 & ~n9436 ;
  assign n11064 = n11062 & n11063 ;
  assign n11065 = n11064 ^ x354 ;
  assign n11066 = n11064 ^ n11062 ;
  assign n11067 = n7474 ^ x1045 ;
  assign n11070 = ~x199 & n11067 ;
  assign n11071 = n11070 ^ x1045 ;
  assign n11072 = n9443 & ~n11071 ;
  assign n11073 = n11072 ^ n3209 ;
  assign n11074 = n11066 & n11073 ;
  assign n11075 = n9441 & n11074 ;
  assign n11076 = n11065 & n11075 ;
  assign n11077 = n11076 ^ n11074 ;
  assign n11078 = n11077 ^ n11073 ;
  assign n11079 = ~n11055 & ~n11078 ;
  assign n11080 = x1111 ^ x723 ;
  assign n11083 = n9162 & ~n11080 ;
  assign n11084 = n11083 ^ x723 ;
  assign n11085 = ~x962 & ~n11084 ;
  assign n11086 = x1114 ^ x724 ;
  assign n11089 = n9162 & ~n11086 ;
  assign n11090 = n11089 ^ x724 ;
  assign n11091 = ~x962 & ~n11090 ;
  assign n11092 = x1120 ^ x725 ;
  assign n11095 = n9162 & ~n11092 ;
  assign n11096 = n11095 ^ x725 ;
  assign n11097 = ~x962 & ~n11096 ;
  assign n11098 = x1126 ^ x726 ;
  assign n11101 = n9162 & n11098 ;
  assign n11102 = n11101 ^ x726 ;
  assign n11103 = ~x962 & n11102 ;
  assign n11104 = x1102 ^ x727 ;
  assign n11107 = n9162 & n11104 ;
  assign n11108 = n11107 ^ x727 ;
  assign n11109 = ~x962 & n11108 ;
  assign n11110 = x1131 ^ x728 ;
  assign n11113 = n9162 & ~n11110 ;
  assign n11114 = n11113 ^ x728 ;
  assign n11115 = ~x962 & ~n11114 ;
  assign n11116 = x1104 ^ x729 ;
  assign n11119 = n9162 & n11116 ;
  assign n11120 = n11119 ^ x729 ;
  assign n11121 = ~x962 & n11120 ;
  assign n11122 = x1106 ^ x730 ;
  assign n11125 = n9162 & n11122 ;
  assign n11126 = n11125 ^ x730 ;
  assign n11127 = ~x962 & n11126 ;
  assign n11128 = ~x945 & x988 ;
  assign n11133 = n11022 & n11128 ;
  assign n11134 = n11133 ^ x731 ;
  assign n11135 = ~n11021 & n11134 ;
  assign n11136 = x1128 ^ x732 ;
  assign n11139 = n9163 & ~n11136 ;
  assign n11140 = n11139 ^ x732 ;
  assign n11141 = ~x962 & ~n11140 ;
  assign n11168 = x399 ^ x375 ;
  assign n11171 = x592 & n11168 ;
  assign n11172 = n11171 ^ x399 ;
  assign n11173 = n9424 & n11172 ;
  assign n11174 = n11173 ^ x316 ;
  assign n11179 = n9441 & n11174 ;
  assign n11175 = x424 & ~n9436 ;
  assign n11177 = n11175 ^ n11173 ;
  assign n11180 = n11179 ^ n11177 ;
  assign n11181 = n11180 ^ x1047 ;
  assign n11165 = x200 & n7845 ;
  assign n11161 = x1047 ^ x308 ;
  assign n11166 = n11165 ^ n11161 ;
  assign n11167 = ~x199 & n11166 ;
  assign n11182 = n11181 ^ n11167 ;
  assign n11183 = ~n9423 & n11182 ;
  assign n11184 = n11183 ^ n11180 ;
  assign n11155 = x838 & n9678 ;
  assign n6101 = x777 ^ x737 ;
  assign n11142 = ~x1135 & n6101 ;
  assign n11143 = n11142 ^ x737 ;
  assign n11145 = n11143 ^ x619 ;
  assign n11144 = n11143 ^ x648 ;
  assign n11146 = n11145 ^ n11144 ;
  assign n11149 = ~x1135 & n11146 ;
  assign n11150 = n11149 ^ n11144 ;
  assign n11151 = ~x1134 & ~n11150 ;
  assign n11152 = n11151 ^ n11143 ;
  assign n11156 = n11155 ^ n11152 ;
  assign n11157 = ~x1136 & ~n11156 ;
  assign n11158 = n11157 ^ n11152 ;
  assign n11159 = n9395 & ~n11158 ;
  assign n11185 = n11184 ^ n11159 ;
  assign n11186 = ~n3209 & n11185 ;
  assign n11187 = n11186 ^ n11184 ;
  assign n11188 = x1119 ^ x734 ;
  assign n11191 = n9162 & ~n11188 ;
  assign n11192 = n11191 ^ x734 ;
  assign n11193 = ~x962 & ~n11192 ;
  assign n11194 = x1109 ^ x735 ;
  assign n11197 = n9162 & n11194 ;
  assign n11198 = n11197 ^ x735 ;
  assign n11199 = ~x962 & n11198 ;
  assign n11200 = x1101 ^ x736 ;
  assign n11203 = n9162 & n11200 ;
  assign n11204 = n11203 ^ x736 ;
  assign n11205 = ~x962 & n11204 ;
  assign n11206 = x1122 ^ x737 ;
  assign n11209 = n9162 & ~n11206 ;
  assign n11210 = n11209 ^ x737 ;
  assign n11211 = ~x962 & ~n11210 ;
  assign n11212 = x1121 ^ x738 ;
  assign n11215 = n9162 & ~n11212 ;
  assign n11216 = n11215 ^ x738 ;
  assign n11217 = ~x962 & ~n11216 ;
  assign n11218 = x1108 ^ x739 ;
  assign n11221 = n8994 & n11218 ;
  assign n11222 = n11221 ^ x739 ;
  assign n11223 = ~x966 & ~n11222 ;
  assign n11224 = x1114 ^ x741 ;
  assign n11227 = n8994 & ~n11224 ;
  assign n11228 = n11227 ^ x741 ;
  assign n11229 = ~x966 & n11228 ;
  assign n11230 = x1112 ^ x742 ;
  assign n11233 = n8994 & ~n11230 ;
  assign n11234 = n11233 ^ x742 ;
  assign n11235 = ~x966 & n11234 ;
  assign n11236 = x1109 ^ x743 ;
  assign n11239 = n8994 & n11236 ;
  assign n11240 = n11239 ^ x743 ;
  assign n11241 = ~x966 & ~n11240 ;
  assign n11242 = x1131 ^ x744 ;
  assign n11245 = n8994 & ~n11242 ;
  assign n11246 = n11245 ^ x744 ;
  assign n11247 = ~x966 & n11246 ;
  assign n11248 = x1111 ^ x745 ;
  assign n11251 = n8994 & ~n11248 ;
  assign n11252 = n11251 ^ x745 ;
  assign n11253 = ~x966 & n11252 ;
  assign n11254 = x1104 ^ x746 ;
  assign n11257 = n8994 & n11254 ;
  assign n11258 = n11257 ^ x746 ;
  assign n11259 = ~x966 & ~n11258 ;
  assign n11264 = x773 & n11128 ;
  assign n11265 = n11264 ^ x747 ;
  assign n11266 = ~n11021 & n11265 ;
  assign n11267 = x1106 ^ x748 ;
  assign n11270 = n8994 & n11267 ;
  assign n11271 = n11270 ^ x748 ;
  assign n11272 = ~x966 & ~n11271 ;
  assign n11273 = x1105 ^ x749 ;
  assign n11276 = n8994 & n11273 ;
  assign n11277 = n11276 ^ x749 ;
  assign n11278 = ~x966 & ~n11277 ;
  assign n11279 = x1130 ^ x750 ;
  assign n11282 = n8994 & ~n11279 ;
  assign n11283 = n11282 ^ x750 ;
  assign n11284 = ~x966 & n11283 ;
  assign n11285 = x1123 ^ x751 ;
  assign n11288 = n8994 & ~n11285 ;
  assign n11289 = n11288 ^ x751 ;
  assign n11290 = ~x966 & n11289 ;
  assign n11291 = x1124 ^ x752 ;
  assign n11294 = n8994 & ~n11291 ;
  assign n11295 = n11294 ^ x752 ;
  assign n11296 = ~x966 & n11295 ;
  assign n11297 = x1117 ^ x753 ;
  assign n11300 = n8994 & ~n11297 ;
  assign n11301 = n11300 ^ x753 ;
  assign n11302 = ~x966 & n11301 ;
  assign n11303 = x1118 ^ x754 ;
  assign n11306 = n8994 & ~n11303 ;
  assign n11307 = n11306 ^ x754 ;
  assign n11308 = ~x966 & n11307 ;
  assign n11309 = x1120 ^ x755 ;
  assign n11312 = n8994 & ~n11309 ;
  assign n11313 = n11312 ^ x755 ;
  assign n11314 = ~x966 & n11313 ;
  assign n11315 = x1119 ^ x756 ;
  assign n11318 = n8994 & ~n11315 ;
  assign n11319 = n11318 ^ x756 ;
  assign n11320 = ~x966 & n11319 ;
  assign n11321 = x1113 ^ x757 ;
  assign n11324 = n8994 & ~n11321 ;
  assign n11325 = n11324 ^ x757 ;
  assign n11326 = ~x966 & n11325 ;
  assign n11327 = x1101 ^ x758 ;
  assign n11330 = n8994 & n11327 ;
  assign n11331 = n11330 ^ x758 ;
  assign n11332 = ~x966 & ~n11331 ;
  assign n11333 = x1100 ^ x759 ;
  assign n11336 = n8994 & n11333 ;
  assign n11337 = n11336 ^ x759 ;
  assign n11338 = ~x966 & ~n11337 ;
  assign n11339 = x1115 ^ x760 ;
  assign n11342 = n8994 & ~n11339 ;
  assign n11343 = n11342 ^ x760 ;
  assign n11344 = ~x966 & n11343 ;
  assign n11345 = x1121 ^ x761 ;
  assign n11348 = n8994 & ~n11345 ;
  assign n11349 = n11348 ^ x761 ;
  assign n11350 = ~x966 & n11349 ;
  assign n11351 = x1129 ^ x762 ;
  assign n11354 = n8994 & ~n11351 ;
  assign n11355 = n11354 ^ x762 ;
  assign n11356 = ~x966 & n11355 ;
  assign n11357 = x1103 ^ x763 ;
  assign n11360 = n8994 & n11357 ;
  assign n11361 = n11360 ^ x763 ;
  assign n11362 = ~x966 & ~n11361 ;
  assign n11363 = x1107 ^ x764 ;
  assign n11366 = n8994 & n11363 ;
  assign n11367 = n11366 ^ x764 ;
  assign n11368 = ~x966 & ~n11367 ;
  assign n11369 = ~x773 & ~x794 ;
  assign n11370 = ~x795 & ~x816 ;
  assign n11371 = n11369 & n11370 ;
  assign n11372 = ~x721 & ~x747 ;
  assign n11374 = x765 & x771 ;
  assign n11373 = x771 ^ x765 ;
  assign n11375 = n11374 ^ n11373 ;
  assign n11376 = n11372 & ~n11375 ;
  assign n11377 = n11371 & n11376 ;
  assign n11378 = n11021 & ~n11377 ;
  assign n11379 = x945 ^ x765 ;
  assign n11380 = ~n11378 & ~n11379 ;
  assign n11381 = x1110 ^ x766 ;
  assign n11384 = n8994 & n11381 ;
  assign n11385 = n11384 ^ x766 ;
  assign n11386 = ~x966 & ~n11385 ;
  assign n11387 = x1116 ^ x767 ;
  assign n11390 = n8994 & ~n11387 ;
  assign n11391 = n11390 ^ x767 ;
  assign n11392 = ~x966 & n11391 ;
  assign n11393 = x1125 ^ x768 ;
  assign n11396 = n8994 & ~n11393 ;
  assign n11397 = n11396 ^ x768 ;
  assign n11398 = ~x966 & n11397 ;
  assign n11399 = n11026 ^ x769 ;
  assign n11400 = ~n11021 & n11399 ;
  assign n11401 = x1126 ^ x770 ;
  assign n11404 = n8994 & ~n11401 ;
  assign n11405 = n11404 ^ x770 ;
  assign n11406 = ~x966 & n11405 ;
  assign n11407 = x987 ^ x771 ;
  assign n11408 = ~x945 & n11407 ;
  assign n11409 = n11408 ^ x771 ;
  assign n11410 = ~n11378 & n11409 ;
  assign n11411 = x1102 ^ x772 ;
  assign n11414 = n8994 & n11411 ;
  assign n11415 = n11414 ^ x772 ;
  assign n11416 = ~x966 & ~n11415 ;
  assign n11417 = n11128 ^ x773 ;
  assign n11418 = ~n11378 & n11417 ;
  assign n11419 = x1127 ^ x774 ;
  assign n11422 = n8994 & ~n11419 ;
  assign n11423 = n11422 ^ x774 ;
  assign n11424 = ~x966 & n11423 ;
  assign n11429 = n11024 & n11374 ;
  assign n11430 = n11429 ^ x775 ;
  assign n11431 = ~n11021 & n11430 ;
  assign n11432 = x1128 ^ x776 ;
  assign n11435 = n8994 & ~n11432 ;
  assign n11436 = n11435 ^ x776 ;
  assign n11437 = ~x966 & n11436 ;
  assign n11438 = x1122 ^ x777 ;
  assign n11441 = n8994 & ~n11438 ;
  assign n11442 = n11441 ^ x777 ;
  assign n11443 = ~x966 & n11442 ;
  assign n11444 = x1100 ^ x778 ;
  assign n11445 = x832 & x956 ;
  assign n11446 = ~x1083 & x1085 ;
  assign n11447 = n11445 & n11446 ;
  assign n11448 = ~x1046 & n11447 ;
  assign n11449 = x968 & n11448 ;
  assign n11450 = n11449 ^ n11448 ;
  assign n11451 = n11444 & n11450 ;
  assign n11452 = n11451 ^ x778 ;
  assign n11453 = x779 & ~n9083 ;
  assign n11454 = x780 & ~n8967 ;
  assign n11455 = x1101 ^ x781 ;
  assign n11456 = n11450 & n11455 ;
  assign n11457 = n11456 ^ x781 ;
  assign n11458 = ~n2649 & ~n8966 ;
  assign n11459 = ~n9010 & n11458 ;
  assign n11460 = x1109 ^ x783 ;
  assign n11461 = n11450 & n11460 ;
  assign n11462 = n11461 ^ x783 ;
  assign n11463 = x1110 ^ x784 ;
  assign n11464 = n11450 & n11463 ;
  assign n11465 = n11464 ^ x784 ;
  assign n11466 = x1102 ^ x785 ;
  assign n11467 = n11450 & n11466 ;
  assign n11468 = n11467 ^ x785 ;
  assign n11469 = x786 ^ x24 ;
  assign n11470 = x954 & n11469 ;
  assign n11471 = n11470 ^ x24 ;
  assign n11472 = x1104 ^ x787 ;
  assign n11473 = n11450 & n11472 ;
  assign n11474 = n11473 ^ x787 ;
  assign n11475 = x1105 ^ x788 ;
  assign n11476 = n11450 & n11475 ;
  assign n11477 = n11476 ^ x788 ;
  assign n11478 = x1106 ^ x789 ;
  assign n11479 = n11450 & n11478 ;
  assign n11480 = n11479 ^ x789 ;
  assign n11481 = x1107 ^ x790 ;
  assign n11482 = n11450 & n11481 ;
  assign n11483 = n11482 ^ x790 ;
  assign n11484 = x1108 ^ x791 ;
  assign n11485 = n11450 & n11484 ;
  assign n11486 = n11485 ^ x791 ;
  assign n11487 = x1103 ^ x792 ;
  assign n11488 = n11450 & n11487 ;
  assign n11489 = n11488 ^ x792 ;
  assign n11490 = x1130 ^ x794 ;
  assign n11491 = n11449 & n11490 ;
  assign n11492 = n11491 ^ x794 ;
  assign n11493 = x1128 ^ x795 ;
  assign n11494 = n11449 & n11493 ;
  assign n11495 = n11494 ^ x795 ;
  assign n11496 = x266 & ~x269 ;
  assign n11497 = x279 & n11496 ;
  assign n11498 = x278 & ~x280 ;
  assign n11499 = n11497 & n11498 ;
  assign n11500 = n9370 & n9372 ;
  assign n11501 = n11499 & n11500 ;
  assign n11502 = n11501 ^ x264 ;
  assign n11503 = x1124 ^ x798 ;
  assign n11504 = n11449 & n11503 ;
  assign n11505 = n11504 ^ x798 ;
  assign n11506 = x1107 ^ x799 ;
  assign n11507 = n11449 & ~n11506 ;
  assign n11508 = n11507 ^ x799 ;
  assign n11509 = x1125 ^ x800 ;
  assign n11510 = n11449 & n11509 ;
  assign n11511 = n11510 ^ x800 ;
  assign n11512 = x1126 ^ x801 ;
  assign n11513 = n11449 & n11512 ;
  assign n11514 = n11513 ^ x801 ;
  assign n11515 = ~x274 & n9375 ;
  assign n11516 = x1106 ^ x803 ;
  assign n11517 = n11449 & ~n11516 ;
  assign n11518 = n11517 ^ x803 ;
  assign n11519 = x1109 ^ x804 ;
  assign n11520 = n11449 & n11519 ;
  assign n11521 = n11520 ^ x804 ;
  assign n11522 = n9371 ^ x270 ;
  assign n11523 = x1127 ^ x807 ;
  assign n11524 = n11449 & n11523 ;
  assign n11525 = n11524 ^ x807 ;
  assign n11526 = x1101 ^ x808 ;
  assign n11527 = n11449 & n11526 ;
  assign n11528 = n11527 ^ x808 ;
  assign n11529 = x1103 ^ x809 ;
  assign n11530 = n11449 & ~n11529 ;
  assign n11531 = n11530 ^ x809 ;
  assign n11532 = x1108 ^ x810 ;
  assign n11533 = n11449 & n11532 ;
  assign n11534 = n11533 ^ x810 ;
  assign n11535 = x1102 ^ x811 ;
  assign n11536 = n11449 & n11535 ;
  assign n11537 = n11536 ^ x811 ;
  assign n11538 = x1104 ^ x812 ;
  assign n11539 = n11449 & ~n11538 ;
  assign n11540 = n11539 ^ x812 ;
  assign n11541 = x1131 ^ x813 ;
  assign n11542 = n11449 & n11541 ;
  assign n11543 = n11542 ^ x813 ;
  assign n11544 = x1105 ^ x814 ;
  assign n11545 = n11449 & ~n11544 ;
  assign n11546 = n11545 ^ x814 ;
  assign n11547 = x1110 ^ x815 ;
  assign n11548 = n11449 & n11547 ;
  assign n11549 = n11548 ^ x815 ;
  assign n11550 = x1129 ^ x816 ;
  assign n11551 = n11449 & n11550 ;
  assign n11552 = n11551 ^ x816 ;
  assign n11553 = n9368 ^ x269 ;
  assign n11554 = n9374 ^ x265 ;
  assign n11555 = ~x270 & n9371 ;
  assign n11556 = n11555 ^ x277 ;
  assign n11557 = ~x811 & ~x893 ;
  assign n11558 = n1844 & n1847 ;
  assign n11559 = n3209 & n11558 ;
  assign n11560 = n11559 ^ n1844 ;
  assign n11562 = ~x982 & ~n1849 ;
  assign n11563 = n11560 & n11562 ;
  assign n11564 = n11563 ^ n11559 ;
  assign n11569 = x1131 ^ x1130 ;
  assign n11568 = x1129 ^ x1128 ;
  assign n11570 = n11569 ^ n11568 ;
  assign n11566 = x1125 ^ x1124 ;
  assign n11565 = x1127 ^ x1126 ;
  assign n11567 = n11566 ^ n11565 ;
  assign n11571 = n11570 ^ n11567 ;
  assign n11572 = n11571 ^ x825 ;
  assign n11573 = x123 & ~x222 ;
  assign n11574 = n9423 & n11573 ;
  assign n11575 = ~n11572 & ~n11574 ;
  assign n11576 = n11575 ^ x825 ;
  assign n11581 = x1123 ^ x1122 ;
  assign n11580 = x1121 ^ x1120 ;
  assign n11582 = n11581 ^ n11580 ;
  assign n11578 = x1117 ^ x1116 ;
  assign n11577 = x1119 ^ x1118 ;
  assign n11579 = n11578 ^ n11577 ;
  assign n11583 = n11582 ^ n11579 ;
  assign n11584 = n11583 ^ x826 ;
  assign n11585 = ~n11574 & ~n11584 ;
  assign n11586 = n11585 ^ x826 ;
  assign n11591 = x1107 ^ x1106 ;
  assign n11590 = x1105 ^ x1104 ;
  assign n11592 = n11591 ^ n11590 ;
  assign n11588 = x1103 ^ x1102 ;
  assign n11587 = x1101 ^ x1100 ;
  assign n11589 = n11588 ^ n11587 ;
  assign n11593 = n11592 ^ n11589 ;
  assign n11594 = n11593 ^ x827 ;
  assign n11595 = ~n11574 & ~n11594 ;
  assign n11596 = n11595 ^ x827 ;
  assign n11601 = x1109 ^ x1108 ;
  assign n11600 = x1111 ^ x1110 ;
  assign n11602 = n11601 ^ n11600 ;
  assign n11598 = x1113 ^ x1112 ;
  assign n11597 = x1115 ^ x1114 ;
  assign n11599 = n11598 ^ n11597 ;
  assign n11603 = n11602 ^ n11599 ;
  assign n11604 = n11603 ^ x828 ;
  assign n11605 = ~n11574 & ~n11604 ;
  assign n11606 = n11605 ^ x828 ;
  assign n11607 = n3209 & n7928 ;
  assign n11608 = ~x951 & x1092 ;
  assign n11609 = ~n11607 & n11608 ;
  assign n11610 = n11609 ^ n11607 ;
  assign n11611 = n11499 ^ x281 ;
  assign n11612 = ~x832 & ~x1163 ;
  assign n11613 = n3010 & n7928 ;
  assign n11614 = n11612 & n11613 ;
  assign n11615 = x1091 ^ x833 ;
  assign n11616 = n3009 & n11615 ;
  assign n11617 = n11616 ^ x833 ;
  assign n11618 = x946 & n3009 ;
  assign n11619 = ~x281 & n9369 ;
  assign n11620 = n11619 ^ x282 ;
  assign n11621 = x1049 ^ x837 ;
  assign n11622 = ~x955 & n11621 ;
  assign n11623 = n11622 ^ x837 ;
  assign n11624 = x1047 ^ x838 ;
  assign n11625 = ~x955 & n11624 ;
  assign n11626 = n11625 ^ x838 ;
  assign n11627 = x1074 ^ x839 ;
  assign n11628 = ~x955 & n11627 ;
  assign n11629 = n11628 ^ x839 ;
  assign n11630 = x1196 ^ x840 ;
  assign n11631 = n3009 & n11630 ;
  assign n11632 = n11631 ^ x840 ;
  assign n11633 = n3543 & n5634 ;
  assign n11634 = x1035 ^ x842 ;
  assign n11635 = ~x955 & n11634 ;
  assign n11636 = n11635 ^ x842 ;
  assign n11637 = x1079 ^ x843 ;
  assign n11638 = ~x955 & n11637 ;
  assign n11639 = n11638 ^ x843 ;
  assign n11640 = x1078 ^ x844 ;
  assign n11641 = ~x955 & n11640 ;
  assign n11642 = n11641 ^ x844 ;
  assign n11643 = x1043 ^ x845 ;
  assign n11644 = ~x955 & n11643 ;
  assign n11645 = n11644 ^ x845 ;
  assign n11646 = x1134 ^ x846 ;
  assign n11647 = ~n7492 & n11646 ;
  assign n11648 = n11647 ^ x846 ;
  assign n11649 = x1055 ^ x847 ;
  assign n11650 = ~x955 & n11649 ;
  assign n11651 = n11650 ^ x847 ;
  assign n11652 = x1039 ^ x848 ;
  assign n11653 = ~x955 & n11652 ;
  assign n11654 = n11653 ^ x848 ;
  assign n11655 = x1198 ^ x849 ;
  assign n11656 = n3009 & n11655 ;
  assign n11657 = n11656 ^ x849 ;
  assign n11658 = x1048 ^ x850 ;
  assign n11659 = ~x955 & n11658 ;
  assign n11660 = n11659 ^ x850 ;
  assign n11661 = x1045 ^ x851 ;
  assign n11662 = ~x955 & n11661 ;
  assign n11663 = n11662 ^ x851 ;
  assign n11664 = x1062 ^ x852 ;
  assign n11665 = ~x955 & n11664 ;
  assign n11666 = n11665 ^ x852 ;
  assign n11667 = x1080 ^ x853 ;
  assign n11668 = ~x955 & n11667 ;
  assign n11669 = n11668 ^ x853 ;
  assign n11670 = x1051 ^ x854 ;
  assign n11671 = ~x955 & n11670 ;
  assign n11672 = n11671 ^ x854 ;
  assign n11673 = x1065 ^ x855 ;
  assign n11674 = ~x955 & n11673 ;
  assign n11675 = n11674 ^ x855 ;
  assign n11676 = x1067 ^ x856 ;
  assign n11677 = ~x955 & n11676 ;
  assign n11678 = n11677 ^ x856 ;
  assign n11679 = x1058 ^ x857 ;
  assign n11680 = ~x955 & n11679 ;
  assign n11681 = n11680 ^ x857 ;
  assign n11682 = x1087 ^ x858 ;
  assign n11683 = ~x955 & n11682 ;
  assign n11684 = n11683 ^ x858 ;
  assign n11685 = x1070 ^ x859 ;
  assign n11686 = ~x955 & n11685 ;
  assign n11687 = n11686 ^ x859 ;
  assign n11688 = x1076 ^ x860 ;
  assign n11689 = ~x955 & n11688 ;
  assign n11690 = n11689 ^ x860 ;
  assign n11691 = x1141 ^ x861 ;
  assign n11692 = ~n7492 & n11691 ;
  assign n11693 = n11692 ^ x861 ;
  assign n11694 = x1139 ^ x862 ;
  assign n11695 = ~n7492 & n11694 ;
  assign n11696 = n11695 ^ x862 ;
  assign n11697 = x1199 ^ x863 ;
  assign n11698 = n3009 & n11697 ;
  assign n11699 = n11698 ^ x863 ;
  assign n11700 = x1197 ^ x864 ;
  assign n11701 = n3009 & n11700 ;
  assign n11702 = n11701 ^ x864 ;
  assign n11703 = x1040 ^ x865 ;
  assign n11704 = ~x955 & n11703 ;
  assign n11705 = n11704 ^ x865 ;
  assign n11706 = x1053 ^ x866 ;
  assign n11707 = ~x955 & n11706 ;
  assign n11708 = n11707 ^ x866 ;
  assign n11709 = x1057 ^ x867 ;
  assign n11710 = ~x955 & n11709 ;
  assign n11711 = n11710 ^ x867 ;
  assign n11712 = x1063 ^ x868 ;
  assign n11713 = ~x955 & n11712 ;
  assign n11714 = n11713 ^ x868 ;
  assign n11715 = x1140 ^ x869 ;
  assign n11716 = ~n7492 & n11715 ;
  assign n11717 = n11716 ^ x869 ;
  assign n11718 = x1069 ^ x870 ;
  assign n11719 = ~x955 & n11718 ;
  assign n11720 = n11719 ^ x870 ;
  assign n11721 = x1072 ^ x871 ;
  assign n11722 = ~x955 & n11721 ;
  assign n11723 = n11722 ^ x871 ;
  assign n11724 = x1084 ^ x872 ;
  assign n11725 = ~x955 & n11724 ;
  assign n11726 = n11725 ^ x872 ;
  assign n11727 = x1044 ^ x873 ;
  assign n11728 = ~x955 & n11727 ;
  assign n11729 = n11728 ^ x873 ;
  assign n11730 = x1036 ^ x874 ;
  assign n11731 = ~x955 & n11730 ;
  assign n11732 = n11731 ^ x874 ;
  assign n11733 = x1136 ^ x875 ;
  assign n11734 = ~n7492 & n11733 ;
  assign n11735 = n11734 ^ x875 ;
  assign n11736 = x1037 ^ x876 ;
  assign n11737 = ~x955 & n11736 ;
  assign n11738 = n11737 ^ x876 ;
  assign n11739 = x1138 ^ x877 ;
  assign n11740 = ~n7492 & n11739 ;
  assign n11741 = n11740 ^ x877 ;
  assign n11742 = x1137 ^ x878 ;
  assign n11743 = ~n7492 & n11742 ;
  assign n11744 = n11743 ^ x878 ;
  assign n11745 = x1135 ^ x879 ;
  assign n11746 = ~n7492 & n11745 ;
  assign n11747 = n11746 ^ x879 ;
  assign n11748 = x1081 ^ x880 ;
  assign n11749 = ~x955 & n11748 ;
  assign n11750 = n11749 ^ x880 ;
  assign n11751 = x1059 ^ x881 ;
  assign n11752 = ~x955 & n11751 ;
  assign n11753 = n11752 ^ x881 ;
  assign n11754 = x1107 ^ x883 ;
  assign n11755 = ~n11574 & ~n11754 ;
  assign n11756 = n11755 ^ x883 ;
  assign n11757 = x1124 ^ x884 ;
  assign n11758 = ~n11574 & ~n11757 ;
  assign n11759 = n11758 ^ x884 ;
  assign n11760 = x1125 ^ x885 ;
  assign n11761 = ~n11574 & ~n11760 ;
  assign n11762 = n11761 ^ x885 ;
  assign n11763 = x1109 ^ x886 ;
  assign n11764 = ~n11574 & ~n11763 ;
  assign n11765 = n11764 ^ x886 ;
  assign n11766 = x1100 ^ x887 ;
  assign n11767 = ~n11574 & ~n11766 ;
  assign n11768 = n11767 ^ x887 ;
  assign n11769 = x1120 ^ x888 ;
  assign n11770 = ~n11574 & ~n11769 ;
  assign n11771 = n11770 ^ x888 ;
  assign n11772 = x1103 ^ x889 ;
  assign n11773 = ~n11574 & ~n11772 ;
  assign n11774 = n11773 ^ x889 ;
  assign n11775 = x1126 ^ x890 ;
  assign n11776 = ~n11574 & ~n11775 ;
  assign n11777 = n11776 ^ x890 ;
  assign n11778 = x1116 ^ x891 ;
  assign n11779 = ~n11574 & ~n11778 ;
  assign n11780 = n11779 ^ x891 ;
  assign n11781 = x1101 ^ x892 ;
  assign n11782 = ~n11574 & ~n11781 ;
  assign n11783 = n11782 ^ x892 ;
  assign n11784 = x1119 ^ x894 ;
  assign n11785 = ~n11574 & ~n11784 ;
  assign n11786 = n11785 ^ x894 ;
  assign n11787 = x1113 ^ x895 ;
  assign n11788 = ~n11574 & ~n11787 ;
  assign n11789 = n11788 ^ x895 ;
  assign n11790 = x1118 ^ x896 ;
  assign n11791 = ~n11574 & ~n11790 ;
  assign n11792 = n11791 ^ x896 ;
  assign n11793 = x1129 ^ x898 ;
  assign n11794 = ~n11574 & ~n11793 ;
  assign n11795 = n11794 ^ x898 ;
  assign n11796 = x1115 ^ x899 ;
  assign n11797 = ~n11574 & ~n11796 ;
  assign n11798 = n11797 ^ x899 ;
  assign n11799 = x1110 ^ x900 ;
  assign n11800 = ~n11574 & ~n11799 ;
  assign n11801 = n11800 ^ x900 ;
  assign n11802 = x1111 ^ x902 ;
  assign n11803 = ~n11574 & ~n11802 ;
  assign n11804 = n11803 ^ x902 ;
  assign n11805 = x1121 ^ x903 ;
  assign n11806 = ~n11574 & ~n11805 ;
  assign n11807 = n11806 ^ x903 ;
  assign n11808 = x1127 ^ x904 ;
  assign n11809 = ~n11574 & ~n11808 ;
  assign n11810 = n11809 ^ x904 ;
  assign n11811 = x1131 ^ x905 ;
  assign n11812 = ~n11574 & ~n11811 ;
  assign n11813 = n11812 ^ x905 ;
  assign n11814 = x1128 ^ x906 ;
  assign n11815 = ~n11574 & ~n11814 ;
  assign n11816 = n11815 ^ x906 ;
  assign n11819 = ~x598 & x979 ;
  assign n11820 = ~x615 & n11819 ;
  assign n11817 = ~x624 & ~x979 ;
  assign n11818 = x604 & n11817 ;
  assign n11821 = n11820 ^ n11818 ;
  assign n11822 = n11821 ^ x907 ;
  assign n11823 = x782 & n11822 ;
  assign n11824 = n11823 ^ x907 ;
  assign n11825 = x1122 ^ x908 ;
  assign n11826 = ~n11574 & ~n11825 ;
  assign n11827 = n11826 ^ x908 ;
  assign n11828 = x1105 ^ x909 ;
  assign n11829 = ~n11574 & ~n11828 ;
  assign n11830 = n11829 ^ x909 ;
  assign n11831 = x1117 ^ x910 ;
  assign n11832 = ~n11574 & ~n11831 ;
  assign n11833 = n11832 ^ x910 ;
  assign n11834 = x1130 ^ x911 ;
  assign n11835 = ~n11574 & ~n11834 ;
  assign n11836 = n11835 ^ x911 ;
  assign n11837 = x1114 ^ x912 ;
  assign n11838 = ~n11574 & ~n11837 ;
  assign n11839 = n11838 ^ x912 ;
  assign n11840 = x1106 ^ x913 ;
  assign n11841 = ~n11574 & ~n11840 ;
  assign n11842 = n11841 ^ x913 ;
  assign n11843 = n9367 ^ x280 ;
  assign n11844 = x1108 ^ x915 ;
  assign n11845 = ~n11574 & ~n11844 ;
  assign n11846 = n11845 ^ x915 ;
  assign n11847 = x1123 ^ x916 ;
  assign n11848 = ~n11574 & ~n11847 ;
  assign n11849 = n11848 ^ x916 ;
  assign n11850 = x1112 ^ x917 ;
  assign n11851 = ~n11574 & ~n11850 ;
  assign n11852 = n11851 ^ x917 ;
  assign n11853 = x1104 ^ x918 ;
  assign n11854 = ~n11574 & ~n11853 ;
  assign n11855 = n11854 ^ x918 ;
  assign n11856 = x1102 ^ x919 ;
  assign n11857 = ~n11574 & ~n11856 ;
  assign n11858 = n11857 ^ x919 ;
  assign n11859 = x1139 ^ x920 ;
  assign n11860 = x1093 & n11859 ;
  assign n11861 = n11860 ^ x920 ;
  assign n11862 = x1140 ^ x921 ;
  assign n11863 = x1093 & n11862 ;
  assign n11864 = n11863 ^ x921 ;
  assign n11865 = x1152 ^ x922 ;
  assign n11866 = x1093 & n11865 ;
  assign n11867 = n11866 ^ x922 ;
  assign n11868 = x1154 ^ x923 ;
  assign n11869 = x1093 & n11868 ;
  assign n11870 = n11869 ^ x923 ;
  assign n11871 = x311 & n7858 ;
  assign n11872 = x1155 ^ x925 ;
  assign n11873 = x1093 & n11872 ;
  assign n11874 = n11873 ^ x925 ;
  assign n11875 = x1157 ^ x926 ;
  assign n11876 = x1093 & n11875 ;
  assign n11877 = n11876 ^ x926 ;
  assign n11878 = x1145 ^ x927 ;
  assign n11879 = x1093 & n11878 ;
  assign n11880 = n11879 ^ x927 ;
  assign n11881 = x1136 ^ x928 ;
  assign n11882 = x1093 & n11881 ;
  assign n11883 = n11882 ^ x928 ;
  assign n11884 = x1144 ^ x929 ;
  assign n11885 = x1093 & n11884 ;
  assign n11886 = n11885 ^ x929 ;
  assign n11887 = x1134 ^ x930 ;
  assign n11888 = x1093 & n11887 ;
  assign n11889 = n11888 ^ x930 ;
  assign n11890 = x1150 ^ x931 ;
  assign n11891 = x1093 & n11890 ;
  assign n11892 = n11891 ^ x931 ;
  assign n11893 = x1093 & n2061 ;
  assign n11894 = n11893 ^ x932 ;
  assign n11895 = x1137 ^ x933 ;
  assign n11896 = x1093 & n11895 ;
  assign n11897 = n11896 ^ x933 ;
  assign n11898 = x1147 ^ x934 ;
  assign n11899 = x1093 & n11898 ;
  assign n11900 = n11899 ^ x934 ;
  assign n11901 = x1141 ^ x935 ;
  assign n11902 = x1093 & n11901 ;
  assign n11903 = n11902 ^ x935 ;
  assign n11904 = x1149 ^ x936 ;
  assign n11905 = x1093 & n11904 ;
  assign n11906 = n11905 ^ x936 ;
  assign n11907 = x1148 ^ x937 ;
  assign n11908 = x1093 & n11907 ;
  assign n11909 = n11908 ^ x937 ;
  assign n11910 = x1135 ^ x938 ;
  assign n11911 = x1093 & n11910 ;
  assign n11912 = n11911 ^ x938 ;
  assign n11913 = x1146 ^ x939 ;
  assign n11914 = x1093 & n11913 ;
  assign n11915 = n11914 ^ x939 ;
  assign n11916 = x1138 ^ x940 ;
  assign n11917 = x1093 & n11916 ;
  assign n11918 = n11917 ^ x940 ;
  assign n11919 = x1153 ^ x941 ;
  assign n11920 = x1093 & n11919 ;
  assign n11921 = n11920 ^ x941 ;
  assign n11922 = x1156 ^ x942 ;
  assign n11923 = x1093 & n11922 ;
  assign n11924 = n11923 ^ x942 ;
  assign n11925 = x1151 ^ x943 ;
  assign n11926 = x1093 & n11925 ;
  assign n11927 = n11926 ^ x943 ;
  assign n11928 = x1143 ^ x944 ;
  assign n11929 = x1093 & n11928 ;
  assign n11930 = n11929 ^ x944 ;
  assign n11931 = x230 & n3009 ;
  assign n11932 = n11819 ^ x947 ;
  assign n11933 = n11932 ^ n11817 ;
  assign n11934 = x782 & ~n11933 ;
  assign n11935 = n11934 ^ x947 ;
  assign n11936 = x992 ^ x266 ;
  assign n11937 = x949 ^ x313 ;
  assign n11938 = x954 & ~n11937 ;
  assign n11939 = n11938 ^ x313 ;
  assign n11940 = x1092 & n1849 ;
  assign n11941 = ~x31 & x957 ;
  assign n11942 = x1092 & n11941 ;
  assign n11943 = n11942 ^ x31 ;
  assign n11944 = ~x782 & x960 ;
  assign n11945 = ~x230 & x961 ;
  assign n11946 = ~x782 & x963 ;
  assign n11947 = ~x230 & x967 ;
  assign n11948 = ~x230 & x969 ;
  assign n11949 = ~x782 & x970 ;
  assign n11950 = ~x230 & x971 ;
  assign n11951 = ~x782 & x972 ;
  assign n11952 = ~x230 & x974 ;
  assign n11953 = ~x782 & x975 ;
  assign n11954 = ~x230 & x977 ;
  assign n11955 = ~x782 & x978 ;
  assign n11956 = ~x598 & x615 ;
  assign n11957 = x824 & x1092 ;
  assign n11958 = ~x604 & ~x624 ;
  assign y0 = x668 ;
  assign y1 = x672 ;
  assign y2 = x664 ;
  assign y3 = x667 ;
  assign y4 = x676 ;
  assign y5 = x673 ;
  assign y6 = x675 ;
  assign y7 = x666 ;
  assign y8 = x679 ;
  assign y9 = x674 ;
  assign y10 = x663 ;
  assign y11 = x670 ;
  assign y12 = x677 ;
  assign y13 = x682 ;
  assign y14 = x671 ;
  assign y15 = x678 ;
  assign y16 = x718 ;
  assign y17 = x707 ;
  assign y18 = x708 ;
  assign y19 = x713 ;
  assign y20 = x711 ;
  assign y21 = x716 ;
  assign y22 = x733 ;
  assign y23 = x712 ;
  assign y24 = x689 ;
  assign y25 = x717 ;
  assign y26 = x692 ;
  assign y27 = x719 ;
  assign y28 = x722 ;
  assign y29 = x714 ;
  assign y30 = x720 ;
  assign y31 = x685 ;
  assign y32 = x837 ;
  assign y33 = x850 ;
  assign y34 = x872 ;
  assign y35 = x871 ;
  assign y36 = x881 ;
  assign y37 = x866 ;
  assign y38 = x876 ;
  assign y39 = x873 ;
  assign y40 = x874 ;
  assign y41 = x859 ;
  assign y42 = x855 ;
  assign y43 = x852 ;
  assign y44 = x870 ;
  assign y45 = x848 ;
  assign y46 = x865 ;
  assign y47 = x856 ;
  assign y48 = x853 ;
  assign y49 = x847 ;
  assign y50 = x857 ;
  assign y51 = x854 ;
  assign y52 = x858 ;
  assign y53 = x845 ;
  assign y54 = x838 ;
  assign y55 = x842 ;
  assign y56 = x843 ;
  assign y57 = x839 ;
  assign y58 = x844 ;
  assign y59 = x868 ;
  assign y60 = x851 ;
  assign y61 = x867 ;
  assign y62 = x880 ;
  assign y63 = x860 ;
  assign y64 = x1030 ;
  assign y65 = x1034 ;
  assign y66 = x1015 ;
  assign y67 = x1020 ;
  assign y68 = x1025 ;
  assign y69 = x1005 ;
  assign y70 = x996 ;
  assign y71 = x1012 ;
  assign y72 = x993 ;
  assign y73 = x1016 ;
  assign y74 = x1021 ;
  assign y75 = x1010 ;
  assign y76 = x1027 ;
  assign y77 = x1018 ;
  assign y78 = x1017 ;
  assign y79 = x1024 ;
  assign y80 = x1009 ;
  assign y81 = x1032 ;
  assign y82 = x1003 ;
  assign y83 = x997 ;
  assign y84 = x1013 ;
  assign y85 = x1011 ;
  assign y86 = x1008 ;
  assign y87 = x1019 ;
  assign y88 = x1031 ;
  assign y89 = x1022 ;
  assign y90 = x1000 ;
  assign y91 = x1023 ;
  assign y92 = x1002 ;
  assign y93 = x1026 ;
  assign y94 = x1006 ;
  assign y95 = x998 ;
  assign y96 = x31 ;
  assign y97 = x80 ;
  assign y98 = x893 ;
  assign y99 = x467 ;
  assign y100 = x78 ;
  assign y101 = x112 ;
  assign y102 = x13 ;
  assign y103 = x25 ;
  assign y104 = x226 ;
  assign y105 = x127 ;
  assign y106 = x822 ;
  assign y107 = x808 ;
  assign y108 = x227 ;
  assign y109 = x477 ;
  assign y110 = x834 ;
  assign y111 = x229 ;
  assign y112 = x12 ;
  assign y113 = x11 ;
  assign y114 = x10 ;
  assign y115 = x9 ;
  assign y116 = x8 ;
  assign y117 = x7 ;
  assign y118 = x6 ;
  assign y119 = x5 ;
  assign y120 = x4 ;
  assign y121 = x3 ;
  assign y122 = x0 ;
  assign y123 = x2 ;
  assign y124 = x1 ;
  assign y125 = x310 ;
  assign y126 = x302 ;
  assign y127 = x475 ;
  assign y128 = x474 ;
  assign y129 = x466 ;
  assign y130 = x473 ;
  assign y131 = x471 ;
  assign y132 = x472 ;
  assign y133 = x470 ;
  assign y134 = x469 ;
  assign y135 = x465 ;
  assign y136 = x1028 ;
  assign y137 = x1033 ;
  assign y138 = x995 ;
  assign y139 = x994 ;
  assign y140 = x28 ;
  assign y141 = x27 ;
  assign y142 = x26 ;
  assign y143 = x29 ;
  assign y144 = x15 ;
  assign y145 = x14 ;
  assign y146 = x21 ;
  assign y147 = x20 ;
  assign y148 = x19 ;
  assign y149 = x18 ;
  assign y150 = x17 ;
  assign y151 = x16 ;
  assign y152 = x1096 ;
  assign y153 = ~n1902 ;
  assign y154 = ~n1962 ;
  assign y155 = ~n1990 ;
  assign y156 = n2058 ;
  assign y157 = n2154 ;
  assign y158 = ~n2216 ;
  assign y159 = n2264 ;
  assign y160 = n2329 ;
  assign y161 = ~n2383 ;
  assign y162 = n2442 ;
  assign y163 = n2499 ;
  assign y164 = ~n2551 ;
  assign y165 = n2603 ;
  assign y166 = ~1'b0 ;
  assign y167 = ~n2742 ;
  assign y168 = x228 ;
  assign y169 = x22 ;
  assign y170 = ~x1090 ;
  assign y171 = ~n2876 ;
  assign y172 = n2895 ;
  assign y173 = ~n2900 ;
  assign y174 = ~n2935 ;
  assign y175 = ~n2939 ;
  assign y176 = ~n2943 ;
  assign y177 = ~n2947 ;
  assign y178 = ~n2951 ;
  assign y179 = x1089 ;
  assign y180 = x23 ;
  assign y181 = ~n2742 ;
  assign y182 = ~n2988 ;
  assign y183 = n2996 ;
  assign y184 = ~n3002 ;
  assign y185 = ~n3004 ;
  assign y186 = ~n3006 ;
  assign y187 = ~n3008 ;
  assign y188 = x37 ;
  assign y189 = ~n3454 ;
  assign y190 = ~n3515 ;
  assign y191 = ~n3712 ;
  assign y192 = n3844 ;
  assign y193 = n3925 ;
  assign y194 = n3931 ;
  assign y195 = ~n2985 ;
  assign y196 = ~n3948 ;
  assign y197 = ~n3987 ;
  assign y198 = n3990 ;
  assign y199 = n4061 ;
  assign y200 = n4104 ;
  assign y201 = n4114 ;
  assign y202 = n4124 ;
  assign y203 = n4125 ;
  assign y204 = n4133 ;
  assign y205 = n4147 ;
  assign y206 = n4148 ;
  assign y207 = n4208 ;
  assign y208 = n4232 ;
  assign y209 = n4236 ;
  assign y210 = n4255 ;
  assign y211 = n4263 ;
  assign y212 = n4270 ;
  assign y213 = n4274 ;
  assign y214 = n4285 ;
  assign y215 = n4291 ;
  assign y216 = n4294 ;
  assign y217 = n4298 ;
  assign y218 = ~n4303 ;
  assign y219 = n4305 ;
  assign y220 = n4312 ;
  assign y221 = ~n4316 ;
  assign y222 = n4319 ;
  assign y223 = n4321 ;
  assign y224 = n4328 ;
  assign y225 = n4333 ;
  assign y226 = n4339 ;
  assign y227 = n4344 ;
  assign y228 = ~n4361 ;
  assign y229 = n4376 ;
  assign y230 = ~n4395 ;
  assign y231 = n4404 ;
  assign y232 = n4419 ;
  assign y233 = n4423 ;
  assign y234 = n4448 ;
  assign y235 = n4451 ;
  assign y236 = n4452 ;
  assign y237 = ~n4591 ;
  assign y238 = n4638 ;
  assign y239 = ~n4643 ;
  assign y240 = n4649 ;
  assign y241 = n4655 ;
  assign y242 = n4656 ;
  assign y243 = n4659 ;
  assign y244 = n4660 ;
  assign y245 = n4661 ;
  assign y246 = n4669 ;
  assign y247 = n4674 ;
  assign y248 = n4676 ;
  assign y249 = n4687 ;
  assign y250 = n4694 ;
  assign y251 = n4699 ;
  assign y252 = n4753 ;
  assign y253 = ~n4822 ;
  assign y254 = n4834 ;
  assign y255 = ~n4838 ;
  assign y256 = n4840 ;
  assign y257 = n4854 ;
  assign y258 = n4876 ;
  assign y259 = n4882 ;
  assign y260 = n4883 ;
  assign y261 = n4884 ;
  assign y262 = ~n4889 ;
  assign y263 = x117 ;
  assign y264 = n4890 ;
  assign y265 = n4314 ;
  assign y266 = n4897 ;
  assign y267 = n4898 ;
  assign y268 = ~n4902 ;
  assign y269 = n4906 ;
  assign y270 = ~n4907 ;
  assign y271 = n4914 ;
  assign y272 = n4916 ;
  assign y273 = n4923 ;
  assign y274 = n4925 ;
  assign y275 = ~n2993 ;
  assign y276 = n5064 ;
  assign y277 = n5087 ;
  assign y278 = ~n5101 ;
  assign y279 = n5164 ;
  assign y280 = n5096 ;
  assign y281 = n5187 ;
  assign y282 = ~n5295 ;
  assign y283 = n5362 ;
  assign y284 = n5374 ;
  assign y285 = x131 ;
  assign y286 = ~n5389 ;
  assign y287 = ~n5441 ;
  assign y288 = ~n5084 ;
  assign y289 = n5489 ;
  assign y290 = n5526 ;
  assign y291 = n5560 ;
  assign y292 = n5580 ;
  assign y293 = n5606 ;
  assign y294 = n5614 ;
  assign y295 = ~n5644 ;
  assign y296 = n5650 ;
  assign y297 = ~n5847 ;
  assign y298 = ~n5858 ;
  assign y299 = n5869 ;
  assign y300 = ~n5880 ;
  assign y301 = n5891 ;
  assign y302 = ~n5902 ;
  assign y303 = n5911 ;
  assign y304 = ~n5922 ;
  assign y305 = ~n5931 ;
  assign y306 = n5956 ;
  assign y307 = n5968 ;
  assign y308 = ~n5979 ;
  assign y309 = n5990 ;
  assign y310 = ~n6001 ;
  assign y311 = n6013 ;
  assign y312 = n6025 ;
  assign y313 = n6037 ;
  assign y314 = ~n6048 ;
  assign y315 = n6060 ;
  assign y316 = ~n6071 ;
  assign y317 = ~n6082 ;
  assign y318 = n6091 ;
  assign y319 = ~n6100 ;
  assign y320 = ~n6111 ;
  assign y321 = ~n6122 ;
  assign y322 = n6132 ;
  assign y323 = n6143 ;
  assign y324 = ~n6154 ;
  assign y325 = ~n6165 ;
  assign y326 = ~n6176 ;
  assign y327 = ~n6187 ;
  assign y328 = ~n6198 ;
  assign y329 = ~n6209 ;
  assign y330 = ~n6218 ;
  assign y331 = n6227 ;
  assign y332 = ~n6236 ;
  assign y333 = ~n6245 ;
  assign y334 = ~n6254 ;
  assign y335 = ~n6263 ;
  assign y336 = ~n6272 ;
  assign y337 = ~n6281 ;
  assign y338 = ~n6290 ;
  assign y339 = ~n6299 ;
  assign y340 = ~n6308 ;
  assign y341 = ~n6317 ;
  assign y342 = ~n6326 ;
  assign y343 = ~n6335 ;
  assign y344 = ~n6344 ;
  assign y345 = ~n6353 ;
  assign y346 = n6362 ;
  assign y347 = ~n6371 ;
  assign y348 = ~n6380 ;
  assign y349 = ~n6389 ;
  assign y350 = ~n6398 ;
  assign y351 = ~n6407 ;
  assign y352 = ~n6424 ;
  assign y353 = n6435 ;
  assign y354 = ~n6444 ;
  assign y355 = n6455 ;
  assign y356 = n6466 ;
  assign y357 = n6477 ;
  assign y358 = n6513 ;
  assign y359 = n6522 ;
  assign y360 = n6529 ;
  assign y361 = n6547 ;
  assign y362 = n6552 ;
  assign y363 = n6561 ;
  assign y364 = ~n6572 ;
  assign y365 = ~n6583 ;
  assign y366 = ~n6594 ;
  assign y367 = n6603 ;
  assign y368 = n6612 ;
  assign y369 = n6622 ;
  assign y370 = n6632 ;
  assign y371 = ~n6641 ;
  assign y372 = n6652 ;
  assign y373 = n6663 ;
  assign y374 = ~n6674 ;
  assign y375 = n6679 ;
  assign y376 = n6689 ;
  assign y377 = n6695 ;
  assign y378 = n6706 ;
  assign y379 = n6715 ;
  assign y380 = n6724 ;
  assign y381 = n6733 ;
  assign y382 = ~n6756 ;
  assign y383 = n6767 ;
  assign y384 = n6788 ;
  assign y385 = n6797 ;
  assign y386 = x232 ;
  assign y387 = n6801 ;
  assign y388 = x236 ;
  assign y389 = ~n6871 ;
  assign y390 = ~n6990 ;
  assign y391 = n7045 ;
  assign y392 = n7092 ;
  assign y393 = n6764 ;
  assign y394 = ~n7182 ;
  assign y395 = n7214 ;
  assign y396 = n7233 ;
  assign y397 = n7260 ;
  assign y398 = n7278 ;
  assign y399 = n7296 ;
  assign y400 = ~n7328 ;
  assign y401 = n7336 ;
  assign y402 = n7354 ;
  assign y403 = n7372 ;
  assign y404 = n7381 ;
  assign y405 = n7399 ;
  assign y406 = n7408 ;
  assign y407 = ~n7411 ;
  assign y408 = n7421 ;
  assign y409 = n7429 ;
  assign y410 = n7438 ;
  assign y411 = n7447 ;
  assign y412 = n7453 ;
  assign y413 = n7459 ;
  assign y414 = n7465 ;
  assign y415 = n7471 ;
  assign y416 = n7477 ;
  assign y417 = n7483 ;
  assign y418 = n7489 ;
  assign y419 = ~n7500 ;
  assign y420 = ~n7509 ;
  assign y421 = ~n7520 ;
  assign y422 = ~n7531 ;
  assign y423 = n7542 ;
  assign y424 = n7551 ;
  assign y425 = n7560 ;
  assign y426 = ~n7571 ;
  assign y427 = ~n7582 ;
  assign y428 = n7591 ;
  assign y429 = n7600 ;
  assign y430 = n7609 ;
  assign y431 = ~n7620 ;
  assign y432 = n7629 ;
  assign y433 = n7638 ;
  assign y434 = ~n7649 ;
  assign y435 = n7660 ;
  assign y436 = n7671 ;
  assign y437 = ~n7682 ;
  assign y438 = ~n7693 ;
  assign y439 = ~n7704 ;
  assign y440 = n7713 ;
  assign y441 = ~n7725 ;
  assign y442 = n7744 ;
  assign y443 = n7751 ;
  assign y444 = n7753 ;
  assign y445 = n7756 ;
  assign y446 = n7764 ;
  assign y447 = n7767 ;
  assign y448 = n7770 ;
  assign y449 = n7773 ;
  assign y450 = n7776 ;
  assign y451 = n7779 ;
  assign y452 = n7782 ;
  assign y453 = n7785 ;
  assign y454 = n7788 ;
  assign y455 = n7791 ;
  assign y456 = ~n7799 ;
  assign y457 = ~n7807 ;
  assign y458 = n7815 ;
  assign y459 = ~n7829 ;
  assign y460 = n7832 ;
  assign y461 = n7835 ;
  assign y462 = n7838 ;
  assign y463 = n7841 ;
  assign y464 = n7844 ;
  assign y465 = n7847 ;
  assign y466 = n7850 ;
  assign y467 = ~n7857 ;
  assign y468 = n7865 ;
  assign y469 = n7867 ;
  assign y470 = ~n7878 ;
  assign y471 = n7879 ;
  assign y472 = n7883 ;
  assign y473 = n7886 ;
  assign y474 = n7890 ;
  assign y475 = n7894 ;
  assign y476 = n7897 ;
  assign y477 = n7900 ;
  assign y478 = n7903 ;
  assign y479 = n7906 ;
  assign y480 = n7909 ;
  assign y481 = n7912 ;
  assign y482 = n7915 ;
  assign y483 = n7918 ;
  assign y484 = n7921 ;
  assign y485 = n7924 ;
  assign y486 = n7927 ;
  assign y487 = n7932 ;
  assign y488 = n7936 ;
  assign y489 = ~n7941 ;
  assign y490 = n7944 ;
  assign y491 = n7947 ;
  assign y492 = n7950 ;
  assign y493 = n7953 ;
  assign y494 = n7956 ;
  assign y495 = n7959 ;
  assign y496 = n7962 ;
  assign y497 = ~n7965 ;
  assign y498 = n7968 ;
  assign y499 = n7971 ;
  assign y500 = n7974 ;
  assign y501 = n7977 ;
  assign y502 = n7980 ;
  assign y503 = n7983 ;
  assign y504 = n7986 ;
  assign y505 = n7989 ;
  assign y506 = n7992 ;
  assign y507 = n7995 ;
  assign y508 = n7998 ;
  assign y509 = n8001 ;
  assign y510 = n8004 ;
  assign y511 = n8007 ;
  assign y512 = n8010 ;
  assign y513 = n8013 ;
  assign y514 = n8016 ;
  assign y515 = n8019 ;
  assign y516 = n8022 ;
  assign y517 = n8025 ;
  assign y518 = n8028 ;
  assign y519 = n8031 ;
  assign y520 = n8034 ;
  assign y521 = n8037 ;
  assign y522 = n8040 ;
  assign y523 = n8043 ;
  assign y524 = n8046 ;
  assign y525 = n8049 ;
  assign y526 = n8052 ;
  assign y527 = n8055 ;
  assign y528 = n8058 ;
  assign y529 = n8061 ;
  assign y530 = n8064 ;
  assign y531 = n8067 ;
  assign y532 = n8070 ;
  assign y533 = n8073 ;
  assign y534 = n8076 ;
  assign y535 = n8079 ;
  assign y536 = n8082 ;
  assign y537 = n8085 ;
  assign y538 = n8088 ;
  assign y539 = n8091 ;
  assign y540 = n8094 ;
  assign y541 = n8097 ;
  assign y542 = n8100 ;
  assign y543 = n8103 ;
  assign y544 = n8106 ;
  assign y545 = n8109 ;
  assign y546 = n8112 ;
  assign y547 = n8115 ;
  assign y548 = n8118 ;
  assign y549 = n8121 ;
  assign y550 = n8124 ;
  assign y551 = n8127 ;
  assign y552 = n8130 ;
  assign y553 = n8133 ;
  assign y554 = n8136 ;
  assign y555 = n8139 ;
  assign y556 = n8142 ;
  assign y557 = n8145 ;
  assign y558 = n8148 ;
  assign y559 = n8151 ;
  assign y560 = n8154 ;
  assign y561 = n8157 ;
  assign y562 = n8160 ;
  assign y563 = n8163 ;
  assign y564 = n8166 ;
  assign y565 = n8169 ;
  assign y566 = n8172 ;
  assign y567 = n8175 ;
  assign y568 = n8178 ;
  assign y569 = n8181 ;
  assign y570 = n8184 ;
  assign y571 = n8187 ;
  assign y572 = n8190 ;
  assign y573 = n8193 ;
  assign y574 = n8196 ;
  assign y575 = n8199 ;
  assign y576 = n8202 ;
  assign y577 = n8205 ;
  assign y578 = n8208 ;
  assign y579 = n8211 ;
  assign y580 = n8214 ;
  assign y581 = n8217 ;
  assign y582 = n8220 ;
  assign y583 = n8223 ;
  assign y584 = n8226 ;
  assign y585 = n8229 ;
  assign y586 = n8232 ;
  assign y587 = n8235 ;
  assign y588 = n8238 ;
  assign y589 = n8241 ;
  assign y590 = n8244 ;
  assign y591 = n8247 ;
  assign y592 = n8250 ;
  assign y593 = n8253 ;
  assign y594 = n8256 ;
  assign y595 = n8259 ;
  assign y596 = n8262 ;
  assign y597 = n8265 ;
  assign y598 = n8268 ;
  assign y599 = n8271 ;
  assign y600 = n8274 ;
  assign y601 = n8277 ;
  assign y602 = n8280 ;
  assign y603 = n8283 ;
  assign y604 = n8286 ;
  assign y605 = n8289 ;
  assign y606 = n8292 ;
  assign y607 = n8295 ;
  assign y608 = n8298 ;
  assign y609 = n8301 ;
  assign y610 = n8304 ;
  assign y611 = n8307 ;
  assign y612 = n8310 ;
  assign y613 = n8313 ;
  assign y614 = n8361 ;
  assign y615 = n8364 ;
  assign y616 = n8367 ;
  assign y617 = n8370 ;
  assign y618 = n8373 ;
  assign y619 = n8376 ;
  assign y620 = n8379 ;
  assign y621 = n8382 ;
  assign y622 = n8387 ;
  assign y623 = n8392 ;
  assign y624 = n8398 ;
  assign y625 = n8401 ;
  assign y626 = n8406 ;
  assign y627 = n8411 ;
  assign y628 = n8416 ;
  assign y629 = n8421 ;
  assign y630 = n8426 ;
  assign y631 = n8431 ;
  assign y632 = n8436 ;
  assign y633 = n8439 ;
  assign y634 = ~n7875 ;
  assign y635 = n8440 ;
  assign y636 = x583 ;
  assign y637 = n7726 ;
  assign y638 = n8443 ;
  assign y639 = n8446 ;
  assign y640 = n8449 ;
  assign y641 = n8452 ;
  assign y642 = n8455 ;
  assign y643 = n8458 ;
  assign y644 = n8461 ;
  assign y645 = n8464 ;
  assign y646 = n8467 ;
  assign y647 = n8470 ;
  assign y648 = n8473 ;
  assign y649 = n8476 ;
  assign y650 = n8479 ;
  assign y651 = n8482 ;
  assign y652 = n8485 ;
  assign y653 = n8488 ;
  assign y654 = n8491 ;
  assign y655 = n8494 ;
  assign y656 = n8497 ;
  assign y657 = n8500 ;
  assign y658 = n8503 ;
  assign y659 = n8506 ;
  assign y660 = n8509 ;
  assign y661 = n8512 ;
  assign y662 = n8515 ;
  assign y663 = n8518 ;
  assign y664 = n8521 ;
  assign y665 = n8524 ;
  assign y666 = n8527 ;
  assign y667 = n8530 ;
  assign y668 = n8533 ;
  assign y669 = n8536 ;
  assign y670 = n8539 ;
  assign y671 = n8542 ;
  assign y672 = n8545 ;
  assign y673 = n8548 ;
  assign y674 = n8551 ;
  assign y675 = n8554 ;
  assign y676 = n8557 ;
  assign y677 = n8560 ;
  assign y678 = n8563 ;
  assign y679 = n8566 ;
  assign y680 = n8569 ;
  assign y681 = n8572 ;
  assign y682 = n8575 ;
  assign y683 = n8578 ;
  assign y684 = n8581 ;
  assign y685 = n8584 ;
  assign y686 = n8587 ;
  assign y687 = n8590 ;
  assign y688 = n8593 ;
  assign y689 = n8596 ;
  assign y690 = n8599 ;
  assign y691 = n8602 ;
  assign y692 = n8605 ;
  assign y693 = n8608 ;
  assign y694 = n8611 ;
  assign y695 = n8614 ;
  assign y696 = n8617 ;
  assign y697 = n8620 ;
  assign y698 = n8623 ;
  assign y699 = n8626 ;
  assign y700 = n8629 ;
  assign y701 = n8632 ;
  assign y702 = n8635 ;
  assign y703 = n8638 ;
  assign y704 = n8641 ;
  assign y705 = n8644 ;
  assign y706 = n8647 ;
  assign y707 = n8650 ;
  assign y708 = n8653 ;
  assign y709 = n8656 ;
  assign y710 = n8659 ;
  assign y711 = n8662 ;
  assign y712 = n8665 ;
  assign y713 = n8668 ;
  assign y714 = n8671 ;
  assign y715 = n8674 ;
  assign y716 = n8677 ;
  assign y717 = n8680 ;
  assign y718 = n8683 ;
  assign y719 = n8686 ;
  assign y720 = n8689 ;
  assign y721 = n8692 ;
  assign y722 = n8695 ;
  assign y723 = n8698 ;
  assign y724 = n8707 ;
  assign y725 = n8710 ;
  assign y726 = n8713 ;
  assign y727 = n8716 ;
  assign y728 = n8719 ;
  assign y729 = n8722 ;
  assign y730 = n8725 ;
  assign y731 = n8728 ;
  assign y732 = n8731 ;
  assign y733 = n8734 ;
  assign y734 = n8737 ;
  assign y735 = n8740 ;
  assign y736 = n8743 ;
  assign y737 = n8746 ;
  assign y738 = n8749 ;
  assign y739 = n8752 ;
  assign y740 = ~n2608 ;
  assign y741 = n8755 ;
  assign y742 = n8758 ;
  assign y743 = n8761 ;
  assign y744 = n8764 ;
  assign y745 = n8772 ;
  assign y746 = ~n8799 ;
  assign y747 = ~n8805 ;
  assign y748 = n8811 ;
  assign y749 = n8816 ;
  assign y750 = ~n8939 ;
  assign y751 = n8947 ;
  assign y752 = n8958 ;
  assign y753 = n8963 ;
  assign y754 = n8965 ;
  assign y755 = n8972 ;
  assign y756 = n8979 ;
  assign y757 = n8981 ;
  assign y758 = n8985 ;
  assign y759 = n8988 ;
  assign y760 = n9005 ;
  assign y761 = ~n9020 ;
  assign y762 = n9022 ;
  assign y763 = n9031 ;
  assign y764 = n9037 ;
  assign y765 = n9043 ;
  assign y766 = n9049 ;
  assign y767 = n9055 ;
  assign y768 = n9061 ;
  assign y769 = n9067 ;
  assign y770 = n9073 ;
  assign y771 = n9082 ;
  assign y772 = n9088 ;
  assign y773 = n9097 ;
  assign y774 = n9106 ;
  assign y775 = n9112 ;
  assign y776 = n9118 ;
  assign y777 = n9124 ;
  assign y778 = n9130 ;
  assign y779 = n9136 ;
  assign y780 = n9142 ;
  assign y781 = ~n9156 ;
  assign y782 = n9168 ;
  assign y783 = n9174 ;
  assign y784 = n9180 ;
  assign y785 = n9186 ;
  assign y786 = n9192 ;
  assign y787 = n9198 ;
  assign y788 = n9204 ;
  assign y789 = n9210 ;
  assign y790 = n9216 ;
  assign y791 = n9222 ;
  assign y792 = n9228 ;
  assign y793 = n9234 ;
  assign y794 = n9240 ;
  assign y795 = n9246 ;
  assign y796 = n9252 ;
  assign y797 = n9258 ;
  assign y798 = n9264 ;
  assign y799 = n9270 ;
  assign y800 = n9276 ;
  assign y801 = n9282 ;
  assign y802 = n9288 ;
  assign y803 = n9294 ;
  assign y804 = n9300 ;
  assign y805 = n9306 ;
  assign y806 = n9312 ;
  assign y807 = n9318 ;
  assign y808 = n9324 ;
  assign y809 = n9330 ;
  assign y810 = n9336 ;
  assign y811 = n9342 ;
  assign y812 = n9348 ;
  assign y813 = n9354 ;
  assign y814 = n9360 ;
  assign y815 = n9366 ;
  assign y816 = ~n9376 ;
  assign y817 = n9382 ;
  assign y818 = n9388 ;
  assign y819 = n9394 ;
  assign y820 = ~n9456 ;
  assign y821 = ~n9504 ;
  assign y822 = n9510 ;
  assign y823 = ~n9558 ;
  assign y824 = n9608 ;
  assign y825 = n9658 ;
  assign y826 = n9664 ;
  assign y827 = ~n9726 ;
  assign y828 = ~n9768 ;
  assign y829 = n9818 ;
  assign y830 = ~n9866 ;
  assign y831 = n9916 ;
  assign y832 = ~n9964 ;
  assign y833 = n10014 ;
  assign y834 = n10057 ;
  assign y835 = ~n10118 ;
  assign y836 = ~n10167 ;
  assign y837 = n10173 ;
  assign y838 = n10179 ;
  assign y839 = ~n10221 ;
  assign y840 = n1851 ;
  assign y841 = n10227 ;
  assign y842 = ~n10273 ;
  assign y843 = n10279 ;
  assign y844 = n10285 ;
  assign y845 = n10291 ;
  assign y846 = n10337 ;
  assign y847 = n10343 ;
  assign y848 = n10349 ;
  assign y849 = ~n10394 ;
  assign y850 = n10400 ;
  assign y851 = n10406 ;
  assign y852 = n10412 ;
  assign y853 = n10418 ;
  assign y854 = n10424 ;
  assign y855 = n10430 ;
  assign y856 = n10436 ;
  assign y857 = n10442 ;
  assign y858 = n10448 ;
  assign y859 = n10454 ;
  assign y860 = n10460 ;
  assign y861 = n10466 ;
  assign y862 = n10472 ;
  assign y863 = n10478 ;
  assign y864 = ~n10524 ;
  assign y865 = n10570 ;
  assign y866 = n10576 ;
  assign y867 = n10582 ;
  assign y868 = ~n10628 ;
  assign y869 = ~n10674 ;
  assign y870 = ~n10720 ;
  assign y871 = n10767 ;
  assign y872 = n10773 ;
  assign y873 = ~n10825 ;
  assign y874 = n10871 ;
  assign y875 = ~n10913 ;
  assign y876 = n10959 ;
  assign y877 = n11006 ;
  assign y878 = n11033 ;
  assign y879 = ~n11079 ;
  assign y880 = n11085 ;
  assign y881 = n11091 ;
  assign y882 = n11097 ;
  assign y883 = n11103 ;
  assign y884 = n11109 ;
  assign y885 = n11115 ;
  assign y886 = n11121 ;
  assign y887 = n11127 ;
  assign y888 = n11135 ;
  assign y889 = n11141 ;
  assign y890 = n11187 ;
  assign y891 = n11193 ;
  assign y892 = n11199 ;
  assign y893 = n11205 ;
  assign y894 = n11211 ;
  assign y895 = n11217 ;
  assign y896 = ~n11223 ;
  assign y897 = n8995 ;
  assign y898 = ~n11229 ;
  assign y899 = ~n11235 ;
  assign y900 = ~n11241 ;
  assign y901 = ~n11247 ;
  assign y902 = ~n11253 ;
  assign y903 = ~n11259 ;
  assign y904 = n11266 ;
  assign y905 = ~n11272 ;
  assign y906 = ~n11278 ;
  assign y907 = ~n11284 ;
  assign y908 = ~n11290 ;
  assign y909 = ~n11296 ;
  assign y910 = ~n11302 ;
  assign y911 = ~n11308 ;
  assign y912 = ~n11314 ;
  assign y913 = ~n11320 ;
  assign y914 = ~n11326 ;
  assign y915 = ~n11332 ;
  assign y916 = ~n11338 ;
  assign y917 = ~n11344 ;
  assign y918 = ~n11350 ;
  assign y919 = ~n11356 ;
  assign y920 = ~n11362 ;
  assign y921 = ~n11368 ;
  assign y922 = n11380 ;
  assign y923 = ~n11386 ;
  assign y924 = ~n11392 ;
  assign y925 = ~n11398 ;
  assign y926 = n11400 ;
  assign y927 = ~n11406 ;
  assign y928 = n11410 ;
  assign y929 = ~n11416 ;
  assign y930 = n11418 ;
  assign y931 = ~n11424 ;
  assign y932 = n11431 ;
  assign y933 = ~n11437 ;
  assign y934 = ~n11443 ;
  assign y935 = n11452 ;
  assign y936 = ~n11453 ;
  assign y937 = ~n11454 ;
  assign y938 = n11457 ;
  assign y939 = ~n11459 ;
  assign y940 = n11462 ;
  assign y941 = n11465 ;
  assign y942 = n11468 ;
  assign y943 = ~n11471 ;
  assign y944 = n11474 ;
  assign y945 = n11477 ;
  assign y946 = n11480 ;
  assign y947 = n11483 ;
  assign y948 = n11486 ;
  assign y949 = n11489 ;
  assign y950 = n2698 ;
  assign y951 = n11492 ;
  assign y952 = n11495 ;
  assign y953 = ~n11502 ;
  assign y954 = n9163 ;
  assign y955 = n11505 ;
  assign y956 = ~n11508 ;
  assign y957 = n11511 ;
  assign y958 = n11514 ;
  assign y959 = n11515 ;
  assign y960 = ~n11518 ;
  assign y961 = n11521 ;
  assign y962 = ~n11522 ;
  assign y963 = n11378 ;
  assign y964 = n11525 ;
  assign y965 = n11528 ;
  assign y966 = ~n11531 ;
  assign y967 = n11534 ;
  assign y968 = n11537 ;
  assign y969 = ~n11540 ;
  assign y970 = n11543 ;
  assign y971 = ~n11546 ;
  assign y972 = n11549 ;
  assign y973 = n11552 ;
  assign y974 = ~n11553 ;
  assign y975 = ~n5093 ;
  assign y976 = ~n11554 ;
  assign y977 = ~n11556 ;
  assign y978 = n11021 ;
  assign y979 = n11557 ;
  assign y980 = n9162 ;
  assign y981 = n11564 ;
  assign y982 = ~n11576 ;
  assign y983 = ~n11586 ;
  assign y984 = ~n11596 ;
  assign y985 = ~n11606 ;
  assign y986 = n11610 ;
  assign y987 = ~n11611 ;
  assign y988 = n8994 ;
  assign y989 = n11614 ;
  assign y990 = n11617 ;
  assign y991 = n11618 ;
  assign y992 = ~n11620 ;
  assign y993 = n11623 ;
  assign y994 = n11626 ;
  assign y995 = n11629 ;
  assign y996 = n11632 ;
  assign y997 = n11633 ;
  assign y998 = n11636 ;
  assign y999 = n11639 ;
  assign y1000 = n11642 ;
  assign y1001 = n11645 ;
  assign y1002 = n11648 ;
  assign y1003 = n11651 ;
  assign y1004 = n11654 ;
  assign y1005 = n11657 ;
  assign y1006 = n11660 ;
  assign y1007 = n11663 ;
  assign y1008 = n11666 ;
  assign y1009 = n11669 ;
  assign y1010 = n11672 ;
  assign y1011 = n11675 ;
  assign y1012 = n11678 ;
  assign y1013 = n11681 ;
  assign y1014 = n11684 ;
  assign y1015 = n11687 ;
  assign y1016 = n11690 ;
  assign y1017 = n11693 ;
  assign y1018 = n11696 ;
  assign y1019 = n11699 ;
  assign y1020 = n11702 ;
  assign y1021 = n11705 ;
  assign y1022 = n11708 ;
  assign y1023 = n11711 ;
  assign y1024 = n11714 ;
  assign y1025 = n11717 ;
  assign y1026 = n11720 ;
  assign y1027 = n11723 ;
  assign y1028 = n11726 ;
  assign y1029 = n11729 ;
  assign y1030 = n11732 ;
  assign y1031 = n11735 ;
  assign y1032 = n11738 ;
  assign y1033 = n11741 ;
  assign y1034 = n11744 ;
  assign y1035 = n11747 ;
  assign y1036 = n11750 ;
  assign y1037 = n11753 ;
  assign y1038 = ~n1290 ;
  assign y1039 = ~n11756 ;
  assign y1040 = ~n11759 ;
  assign y1041 = ~n11762 ;
  assign y1042 = ~n11765 ;
  assign y1043 = ~n11768 ;
  assign y1044 = ~n11771 ;
  assign y1045 = ~n11774 ;
  assign y1046 = ~n11777 ;
  assign y1047 = ~n11780 ;
  assign y1048 = ~n11783 ;
  assign y1049 = ~n6809 ;
  assign y1050 = ~n11786 ;
  assign y1051 = ~n11789 ;
  assign y1052 = ~n11792 ;
  assign y1053 = x67 ;
  assign y1054 = ~n11795 ;
  assign y1055 = ~n11798 ;
  assign y1056 = ~n11801 ;
  assign y1057 = ~n2619 ;
  assign y1058 = ~n11804 ;
  assign y1059 = ~n11807 ;
  assign y1060 = ~n11810 ;
  assign y1061 = ~n11813 ;
  assign y1062 = ~n11816 ;
  assign y1063 = n11824 ;
  assign y1064 = ~n11827 ;
  assign y1065 = ~n11830 ;
  assign y1066 = ~n11833 ;
  assign y1067 = ~n11836 ;
  assign y1068 = ~n11839 ;
  assign y1069 = ~n11842 ;
  assign y1070 = ~n11843 ;
  assign y1071 = ~n11846 ;
  assign y1072 = ~n11849 ;
  assign y1073 = ~n11852 ;
  assign y1074 = ~n11855 ;
  assign y1075 = ~n11858 ;
  assign y1076 = n11861 ;
  assign y1077 = n11864 ;
  assign y1078 = n11867 ;
  assign y1079 = n11870 ;
  assign y1080 = n11871 ;
  assign y1081 = n11874 ;
  assign y1082 = n11877 ;
  assign y1083 = n11880 ;
  assign y1084 = n11883 ;
  assign y1085 = n11886 ;
  assign y1086 = n11889 ;
  assign y1087 = n11892 ;
  assign y1088 = n11894 ;
  assign y1089 = n11897 ;
  assign y1090 = n11900 ;
  assign y1091 = n11903 ;
  assign y1092 = n11906 ;
  assign y1093 = n11909 ;
  assign y1094 = n11912 ;
  assign y1095 = n11915 ;
  assign y1096 = n11918 ;
  assign y1097 = n11921 ;
  assign y1098 = n11924 ;
  assign y1099 = n11927 ;
  assign y1100 = n11930 ;
  assign y1101 = ~n2669 ;
  assign y1102 = n11931 ;
  assign y1103 = n11935 ;
  assign y1104 = n11936 ;
  assign y1105 = ~n11939 ;
  assign y1106 = n11940 ;
  assign y1107 = n2694 ;
  assign y1108 = x1134 ;
  assign y1109 = x964 ;
  assign y1110 = ~x954 ;
  assign y1111 = x965 ;
  assign y1112 = n11943 ;
  assign y1113 = x991 ;
  assign y1114 = x985 ;
  assign y1115 = n11944 ;
  assign y1116 = n11945 ;
  assign y1117 = x1014 ;
  assign y1118 = n11946 ;
  assign y1119 = x1029 ;
  assign y1120 = x1004 ;
  assign y1121 = x1007 ;
  assign y1122 = n11947 ;
  assign y1123 = x1135 ;
  assign y1124 = n11948 ;
  assign y1125 = n11949 ;
  assign y1126 = n11950 ;
  assign y1127 = n11951 ;
  assign y1128 = n11952 ;
  assign y1129 = n11953 ;
  assign y1130 = ~x278 ;
  assign y1131 = n11954 ;
  assign y1132 = n11955 ;
  assign y1133 = ~n11956 ;
  assign y1134 = x1064 ;
  assign y1135 = n11957 ;
  assign y1136 = x299 ;
  assign y1137 = ~n11958 ;
  assign y1138 = x1075 ;
  assign y1139 = x1052 ;
  assign y1140 = x771 ;
  assign y1141 = x765 ;
  assign y1142 = x605 ;
  assign y1143 = x601 ;
  assign y1144 = x278 ;
  assign y1145 = x279 ;
  assign y1146 = ~x915 ;
  assign y1147 = ~x825 ;
  assign y1148 = ~x826 ;
  assign y1149 = ~x913 ;
  assign y1150 = ~x894 ;
  assign y1151 = ~x905 ;
  assign y1152 = x1095 ;
  assign y1153 = ~x890 ;
  assign y1154 = x1094 ;
  assign y1155 = ~x906 ;
  assign y1156 = ~x896 ;
  assign y1157 = ~x909 ;
  assign y1158 = ~x911 ;
  assign y1159 = ~x908 ;
  assign y1160 = ~x891 ;
  assign y1161 = ~x902 ;
  assign y1162 = ~x903 ;
  assign y1163 = ~x883 ;
  assign y1164 = ~x888 ;
  assign y1165 = ~x919 ;
  assign y1166 = ~x886 ;
  assign y1167 = ~x912 ;
  assign y1168 = ~x895 ;
  assign y1169 = ~x916 ;
  assign y1170 = ~x889 ;
  assign y1171 = ~x900 ;
  assign y1172 = ~x885 ;
  assign y1173 = ~x904 ;
  assign y1174 = ~x899 ;
  assign y1175 = ~x918 ;
  assign y1176 = ~x898 ;
  assign y1177 = ~x917 ;
  assign y1178 = ~x827 ;
  assign y1179 = ~x887 ;
  assign y1180 = ~x884 ;
  assign y1181 = ~x910 ;
  assign y1182 = ~x828 ;
  assign y1183 = ~x892 ;
  assign y1184 = x1187 ;
  assign y1185 = x1172 ;
  assign y1186 = x1170 ;
  assign y1187 = x1138 ;
  assign y1188 = x1177 ;
  assign y1189 = x1178 ;
  assign y1190 = x863 ;
  assign y1191 = x1203 ;
  assign y1192 = x1185 ;
  assign y1193 = x1171 ;
  assign y1194 = x1192 ;
  assign y1195 = x1137 ;
  assign y1196 = x1186 ;
  assign y1197 = x1165 ;
  assign y1198 = x1164 ;
  assign y1199 = x1098 ;
  assign y1200 = x1183 ;
  assign y1201 = x230 ;
  assign y1202 = x1169 ;
  assign y1203 = x1136 ;
  assign y1204 = x1181 ;
  assign y1205 = x849 ;
  assign y1206 = x1193 ;
  assign y1207 = x1182 ;
  assign y1208 = x1168 ;
  assign y1209 = x1175 ;
  assign y1210 = x1191 ;
  assign y1211 = x1099 ;
  assign y1212 = x1174 ;
  assign y1213 = x1179 ;
  assign y1214 = x1202 ;
  assign y1215 = x1176 ;
  assign y1216 = x1173 ;
  assign y1217 = x1201 ;
  assign y1218 = x1167 ;
  assign y1219 = x840 ;
  assign y1220 = x1189 ;
  assign y1221 = x1195 ;
  assign y1222 = x864 ;
  assign y1223 = x1190 ;
  assign y1224 = x1188 ;
  assign y1225 = x1180 ;
  assign y1226 = x1194 ;
  assign y1227 = x1097 ;
  assign y1228 = x1166 ;
  assign y1229 = x1200 ;
  assign y1230 = x1184 ;
endmodule
