module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 ;
  assign n9 = x6 & ~x7 ;
  assign n10 = n9 ^ x7 ;
  assign n11 = n10 ^ x6 ;
  assign n12 = x2 & x3 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n11 & ~n14 ;
  assign n16 = x4 & ~x5 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = x0 & x1 ;
  assign n21 = n20 ^ x1 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n15 & n23 ;
  assign n25 = n11 & ~n19 ;
  assign n26 = n20 ^ x0 ;
  assign n27 = ~n14 & n26 ;
  assign n28 = n25 & n27 ;
  assign n29 = ~n14 & n21 ;
  assign n30 = n25 & n29 ;
  assign n31 = ~n14 & n20 ;
  assign n32 = n25 & n31 ;
  assign n33 = n12 ^ x2 ;
  assign n34 = ~n22 & n33 ;
  assign n35 = n25 & n34 ;
  assign n36 = n26 & n33 ;
  assign n37 = n25 & n36 ;
  assign n38 = n21 & n33 ;
  assign n39 = n25 & n38 ;
  assign n40 = n20 & n33 ;
  assign n41 = n25 & n40 ;
  assign n42 = n13 & ~n22 ;
  assign n43 = n25 & n42 ;
  assign n44 = n13 & n26 ;
  assign n45 = n25 & n44 ;
  assign n46 = n13 & n21 ;
  assign n47 = n25 & n46 ;
  assign n48 = n13 & n20 ;
  assign n49 = n25 & n48 ;
  assign n50 = n12 & ~n22 ;
  assign n51 = n25 & n50 ;
  assign n52 = n12 & n26 ;
  assign n53 = n25 & n52 ;
  assign n54 = n12 & n21 ;
  assign n55 = n25 & n54 ;
  assign n56 = n12 & n20 ;
  assign n57 = n25 & n56 ;
  assign n58 = ~x5 & ~x6 ;
  assign n59 = ~n14 & n58 ;
  assign n60 = x4 & ~x7 ;
  assign n61 = n60 ^ x4 ;
  assign n62 = ~n22 & n61 ;
  assign n63 = n59 & n62 ;
  assign n64 = n26 & n61 ;
  assign n65 = n59 & n64 ;
  assign n66 = n21 & n61 ;
  assign n67 = n59 & n66 ;
  assign n68 = n20 & n61 ;
  assign n69 = n59 & n68 ;
  assign n70 = n33 & n58 ;
  assign n71 = n62 & n70 ;
  assign n72 = n64 & n70 ;
  assign n73 = n66 & n70 ;
  assign n74 = n68 & n70 ;
  assign n75 = n13 & n58 ;
  assign n76 = n62 & n75 ;
  assign n77 = n64 & n75 ;
  assign n78 = n66 & n75 ;
  assign n79 = n68 & n75 ;
  assign n80 = n12 & n58 ;
  assign n81 = n62 & n80 ;
  assign n82 = n64 & n80 ;
  assign n83 = n66 & n80 ;
  assign n84 = n68 & n80 ;
  assign n85 = n18 & ~n22 ;
  assign n86 = n15 & n85 ;
  assign n87 = n11 & n26 ;
  assign n88 = ~n14 & n18 ;
  assign n89 = n87 & n88 ;
  assign n90 = n11 & n21 ;
  assign n91 = n88 & n90 ;
  assign n92 = n11 & n20 ;
  assign n93 = n88 & n92 ;
  assign n94 = n11 & ~n22 ;
  assign n95 = n18 & n33 ;
  assign n96 = n94 & n95 ;
  assign n97 = n87 & n95 ;
  assign n98 = n90 & n95 ;
  assign n99 = n92 & n95 ;
  assign n100 = n13 & n18 ;
  assign n101 = n94 & n100 ;
  assign n102 = n87 & n100 ;
  assign n103 = n90 & n100 ;
  assign n104 = n92 & n100 ;
  assign n105 = n12 & n18 ;
  assign n106 = n94 & n105 ;
  assign n107 = n87 & n105 ;
  assign n108 = n90 & n105 ;
  assign n109 = n92 & n105 ;
  assign n110 = ~n14 & n17 ;
  assign n111 = n94 & n110 ;
  assign n112 = n87 & n110 ;
  assign n113 = n90 & n110 ;
  assign n114 = n92 & n110 ;
  assign n115 = n17 & n33 ;
  assign n116 = n94 & n115 ;
  assign n117 = n87 & n115 ;
  assign n118 = n90 & n115 ;
  assign n119 = n92 & n115 ;
  assign n120 = n13 & n17 ;
  assign n121 = n94 & n120 ;
  assign n122 = n87 & n120 ;
  assign n123 = n90 & n120 ;
  assign n124 = n92 & n120 ;
  assign n125 = n12 & n17 ;
  assign n126 = n94 & n125 ;
  assign n127 = n87 & n125 ;
  assign n128 = n90 & n125 ;
  assign n129 = n92 & n125 ;
  assign n130 = n9 ^ x6 ;
  assign n131 = ~n14 & n130 ;
  assign n132 = n23 & n131 ;
  assign n133 = ~n19 & n26 ;
  assign n134 = n131 & n133 ;
  assign n135 = ~n19 & n21 ;
  assign n136 = n131 & n135 ;
  assign n137 = ~n19 & n20 ;
  assign n138 = n131 & n137 ;
  assign n139 = n33 & n130 ;
  assign n140 = n23 & n139 ;
  assign n141 = n133 & n139 ;
  assign n142 = n135 & n139 ;
  assign n143 = n137 & n139 ;
  assign n144 = n13 & n130 ;
  assign n145 = n23 & n144 ;
  assign n146 = n133 & n144 ;
  assign n147 = n135 & n144 ;
  assign n148 = n137 & n144 ;
  assign n149 = n12 & n130 ;
  assign n150 = n23 & n149 ;
  assign n151 = n133 & n149 ;
  assign n152 = n135 & n149 ;
  assign n153 = n137 & n149 ;
  assign n154 = n16 & ~n22 ;
  assign n155 = n131 & n154 ;
  assign n156 = n16 & n26 ;
  assign n157 = n131 & n156 ;
  assign n158 = n16 & n21 ;
  assign n159 = n131 & n158 ;
  assign n160 = n16 & n20 ;
  assign n161 = n131 & n160 ;
  assign n162 = n139 & n154 ;
  assign n163 = n139 & n156 ;
  assign n164 = n139 & n158 ;
  assign n165 = n139 & n160 ;
  assign n166 = n144 & n154 ;
  assign n167 = n144 & n156 ;
  assign n168 = n144 & n158 ;
  assign n169 = n144 & n160 ;
  assign n170 = n149 & n154 ;
  assign n171 = n149 & n156 ;
  assign n172 = n149 & n158 ;
  assign n173 = n149 & n160 ;
  assign n174 = n85 & n131 ;
  assign n175 = n26 & n130 ;
  assign n176 = n88 & n175 ;
  assign n177 = n21 & n130 ;
  assign n178 = n88 & n177 ;
  assign n179 = n20 & n130 ;
  assign n180 = n88 & n179 ;
  assign n181 = n85 & n139 ;
  assign n182 = n95 & n175 ;
  assign n183 = n95 & n177 ;
  assign n184 = n95 & n179 ;
  assign n185 = n85 & n144 ;
  assign n186 = n100 & n175 ;
  assign n187 = n100 & n177 ;
  assign n188 = n100 & n179 ;
  assign n189 = n85 & n149 ;
  assign n190 = n105 & n175 ;
  assign n191 = n105 & n177 ;
  assign n192 = n105 & n179 ;
  assign n193 = ~n14 & ~n22 ;
  assign n194 = n17 & n130 ;
  assign n195 = n193 & n194 ;
  assign n196 = n27 & n194 ;
  assign n197 = n29 & n194 ;
  assign n198 = n31 & n194 ;
  assign n199 = n34 & n194 ;
  assign n200 = n36 & n194 ;
  assign n201 = n38 & n194 ;
  assign n202 = n115 & n179 ;
  assign n203 = n42 & n194 ;
  assign n204 = n44 & n194 ;
  assign n205 = n120 & n177 ;
  assign n206 = n48 & n194 ;
  assign n207 = n50 & n194 ;
  assign n208 = n52 & n194 ;
  assign n209 = n54 & n194 ;
  assign n210 = n56 & n194 ;
  assign n211 = ~n10 & ~n19 ;
  assign n212 = n193 & n211 ;
  assign n213 = n27 & n211 ;
  assign n214 = n29 & n211 ;
  assign n215 = n31 & n211 ;
  assign n216 = n34 & n211 ;
  assign n217 = n36 & n211 ;
  assign n218 = n38 & n211 ;
  assign n219 = n40 & n211 ;
  assign n220 = n42 & n211 ;
  assign n221 = n44 & n211 ;
  assign n222 = n46 & n211 ;
  assign n223 = n48 & n211 ;
  assign n224 = n50 & n211 ;
  assign n225 = n52 & n211 ;
  assign n226 = n54 & n211 ;
  assign n227 = n56 & n211 ;
  assign n228 = ~n22 & n60 ;
  assign n229 = n59 & n228 ;
  assign n230 = n26 & n60 ;
  assign n231 = n59 & n230 ;
  assign n232 = n21 & n60 ;
  assign n233 = n59 & n232 ;
  assign n234 = n20 & n60 ;
  assign n235 = n59 & n234 ;
  assign n236 = n70 & n228 ;
  assign n237 = n70 & n230 ;
  assign n238 = n70 & n232 ;
  assign n239 = n70 & n234 ;
  assign n240 = n75 & n228 ;
  assign n241 = n75 & n230 ;
  assign n242 = n75 & n232 ;
  assign n243 = n75 & n234 ;
  assign n244 = n80 & n228 ;
  assign n245 = n80 & n230 ;
  assign n246 = n80 & n232 ;
  assign n247 = n80 & n234 ;
  assign n248 = ~n10 & n18 ;
  assign n249 = n193 & n248 ;
  assign n250 = n27 & n248 ;
  assign n251 = n29 & n248 ;
  assign n252 = n31 & n248 ;
  assign n253 = n34 & n248 ;
  assign n254 = n36 & n248 ;
  assign n255 = n38 & n248 ;
  assign n256 = n40 & n248 ;
  assign n257 = n42 & n248 ;
  assign n258 = n44 & n248 ;
  assign n259 = n46 & n248 ;
  assign n260 = n48 & n248 ;
  assign n261 = n50 & n248 ;
  assign n262 = n52 & n248 ;
  assign n263 = n54 & n248 ;
  assign n264 = n56 & n248 ;
  assign n265 = ~n10 & n17 ;
  assign n266 = n193 & n265 ;
  assign n267 = n27 & n265 ;
  assign n268 = n29 & n265 ;
  assign n269 = n31 & n265 ;
  assign n270 = n34 & n265 ;
  assign n271 = n36 & n265 ;
  assign n272 = n38 & n265 ;
  assign n273 = n40 & n265 ;
  assign n274 = n42 & n265 ;
  assign n275 = n44 & n265 ;
  assign n276 = n46 & n265 ;
  assign n277 = n48 & n265 ;
  assign n278 = n50 & n265 ;
  assign n279 = n52 & n265 ;
  assign n280 = n54 & n265 ;
  assign n281 = n56 & n265 ;
  assign n282 = n9 & ~n19 ;
  assign n283 = n193 & n282 ;
  assign n284 = n27 & n282 ;
  assign n285 = n29 & n282 ;
  assign n286 = n31 & n282 ;
  assign n287 = n34 & n282 ;
  assign n288 = n36 & n282 ;
  assign n289 = n38 & n282 ;
  assign n290 = n40 & n282 ;
  assign n291 = n42 & n282 ;
  assign n292 = n44 & n282 ;
  assign n293 = n46 & n282 ;
  assign n294 = n48 & n282 ;
  assign n295 = n50 & n282 ;
  assign n296 = n52 & n282 ;
  assign n297 = n54 & n282 ;
  assign n298 = n56 & n282 ;
  assign n299 = n9 & n16 ;
  assign n300 = n193 & n299 ;
  assign n301 = n27 & n299 ;
  assign n302 = n29 & n299 ;
  assign n303 = n31 & n299 ;
  assign n304 = n34 & n299 ;
  assign n305 = n36 & n299 ;
  assign n306 = n38 & n299 ;
  assign n307 = n40 & n299 ;
  assign n308 = n42 & n299 ;
  assign n309 = n44 & n299 ;
  assign n310 = n46 & n299 ;
  assign n311 = n48 & n299 ;
  assign n312 = n50 & n299 ;
  assign n313 = n52 & n299 ;
  assign n314 = n54 & n299 ;
  assign n315 = n56 & n299 ;
  assign n316 = n9 & n18 ;
  assign n317 = n193 & n316 ;
  assign n318 = n27 & n316 ;
  assign n319 = n29 & n316 ;
  assign n320 = n31 & n316 ;
  assign n321 = n34 & n316 ;
  assign n322 = n36 & n316 ;
  assign n323 = n38 & n316 ;
  assign n324 = n40 & n316 ;
  assign n325 = n42 & n316 ;
  assign n326 = n44 & n316 ;
  assign n327 = n46 & n316 ;
  assign n328 = n48 & n316 ;
  assign n329 = n50 & n316 ;
  assign n330 = n52 & n316 ;
  assign n331 = n54 & n316 ;
  assign n332 = n56 & n316 ;
  assign n333 = n9 & n17 ;
  assign n334 = n193 & n333 ;
  assign n335 = n27 & n333 ;
  assign n336 = n29 & n333 ;
  assign n337 = n31 & n333 ;
  assign n338 = n34 & n333 ;
  assign n339 = n36 & n333 ;
  assign n340 = n38 & n333 ;
  assign n341 = n40 & n333 ;
  assign n342 = n42 & n333 ;
  assign n343 = n44 & n333 ;
  assign n344 = n46 & n333 ;
  assign n345 = n48 & n333 ;
  assign n346 = n50 & n333 ;
  assign n347 = n52 & n333 ;
  assign n348 = n54 & n333 ;
  assign n349 = n56 & n333 ;
  assign y0 = n24 ;
  assign y1 = n28 ;
  assign y2 = n30 ;
  assign y3 = n32 ;
  assign y4 = n35 ;
  assign y5 = n37 ;
  assign y6 = n39 ;
  assign y7 = n41 ;
  assign y8 = n43 ;
  assign y9 = n45 ;
  assign y10 = n47 ;
  assign y11 = n49 ;
  assign y12 = n51 ;
  assign y13 = n53 ;
  assign y14 = n55 ;
  assign y15 = n57 ;
  assign y16 = n63 ;
  assign y17 = n65 ;
  assign y18 = n67 ;
  assign y19 = n69 ;
  assign y20 = n71 ;
  assign y21 = n72 ;
  assign y22 = n73 ;
  assign y23 = n74 ;
  assign y24 = n76 ;
  assign y25 = n77 ;
  assign y26 = n78 ;
  assign y27 = n79 ;
  assign y28 = n81 ;
  assign y29 = n82 ;
  assign y30 = n83 ;
  assign y31 = n84 ;
  assign y32 = n86 ;
  assign y33 = n89 ;
  assign y34 = n91 ;
  assign y35 = n93 ;
  assign y36 = n96 ;
  assign y37 = n97 ;
  assign y38 = n98 ;
  assign y39 = n99 ;
  assign y40 = n101 ;
  assign y41 = n102 ;
  assign y42 = n103 ;
  assign y43 = n104 ;
  assign y44 = n106 ;
  assign y45 = n107 ;
  assign y46 = n108 ;
  assign y47 = n109 ;
  assign y48 = n111 ;
  assign y49 = n112 ;
  assign y50 = n113 ;
  assign y51 = n114 ;
  assign y52 = n116 ;
  assign y53 = n117 ;
  assign y54 = n118 ;
  assign y55 = n119 ;
  assign y56 = n121 ;
  assign y57 = n122 ;
  assign y58 = n123 ;
  assign y59 = n124 ;
  assign y60 = n126 ;
  assign y61 = n127 ;
  assign y62 = n128 ;
  assign y63 = n129 ;
  assign y64 = n132 ;
  assign y65 = n134 ;
  assign y66 = n136 ;
  assign y67 = n138 ;
  assign y68 = n140 ;
  assign y69 = n141 ;
  assign y70 = n142 ;
  assign y71 = n143 ;
  assign y72 = n145 ;
  assign y73 = n146 ;
  assign y74 = n147 ;
  assign y75 = n148 ;
  assign y76 = n150 ;
  assign y77 = n151 ;
  assign y78 = n152 ;
  assign y79 = n153 ;
  assign y80 = n155 ;
  assign y81 = n157 ;
  assign y82 = n159 ;
  assign y83 = n161 ;
  assign y84 = n162 ;
  assign y85 = n163 ;
  assign y86 = n164 ;
  assign y87 = n165 ;
  assign y88 = n166 ;
  assign y89 = n167 ;
  assign y90 = n168 ;
  assign y91 = n169 ;
  assign y92 = n170 ;
  assign y93 = n171 ;
  assign y94 = n172 ;
  assign y95 = n173 ;
  assign y96 = n174 ;
  assign y97 = n176 ;
  assign y98 = n178 ;
  assign y99 = n180 ;
  assign y100 = n181 ;
  assign y101 = n182 ;
  assign y102 = n183 ;
  assign y103 = n184 ;
  assign y104 = n185 ;
  assign y105 = n186 ;
  assign y106 = n187 ;
  assign y107 = n188 ;
  assign y108 = n189 ;
  assign y109 = n190 ;
  assign y110 = n191 ;
  assign y111 = n192 ;
  assign y112 = n195 ;
  assign y113 = n196 ;
  assign y114 = n197 ;
  assign y115 = n198 ;
  assign y116 = n199 ;
  assign y117 = n200 ;
  assign y118 = n201 ;
  assign y119 = n202 ;
  assign y120 = n203 ;
  assign y121 = n204 ;
  assign y122 = n205 ;
  assign y123 = n206 ;
  assign y124 = n207 ;
  assign y125 = n208 ;
  assign y126 = n209 ;
  assign y127 = n210 ;
  assign y128 = n212 ;
  assign y129 = n213 ;
  assign y130 = n214 ;
  assign y131 = n215 ;
  assign y132 = n216 ;
  assign y133 = n217 ;
  assign y134 = n218 ;
  assign y135 = n219 ;
  assign y136 = n220 ;
  assign y137 = n221 ;
  assign y138 = n222 ;
  assign y139 = n223 ;
  assign y140 = n224 ;
  assign y141 = n225 ;
  assign y142 = n226 ;
  assign y143 = n227 ;
  assign y144 = n229 ;
  assign y145 = n231 ;
  assign y146 = n233 ;
  assign y147 = n235 ;
  assign y148 = n236 ;
  assign y149 = n237 ;
  assign y150 = n238 ;
  assign y151 = n239 ;
  assign y152 = n240 ;
  assign y153 = n241 ;
  assign y154 = n242 ;
  assign y155 = n243 ;
  assign y156 = n244 ;
  assign y157 = n245 ;
  assign y158 = n246 ;
  assign y159 = n247 ;
  assign y160 = n249 ;
  assign y161 = n250 ;
  assign y162 = n251 ;
  assign y163 = n252 ;
  assign y164 = n253 ;
  assign y165 = n254 ;
  assign y166 = n255 ;
  assign y167 = n256 ;
  assign y168 = n257 ;
  assign y169 = n258 ;
  assign y170 = n259 ;
  assign y171 = n260 ;
  assign y172 = n261 ;
  assign y173 = n262 ;
  assign y174 = n263 ;
  assign y175 = n264 ;
  assign y176 = n266 ;
  assign y177 = n267 ;
  assign y178 = n268 ;
  assign y179 = n269 ;
  assign y180 = n270 ;
  assign y181 = n271 ;
  assign y182 = n272 ;
  assign y183 = n273 ;
  assign y184 = n274 ;
  assign y185 = n275 ;
  assign y186 = n276 ;
  assign y187 = n277 ;
  assign y188 = n278 ;
  assign y189 = n279 ;
  assign y190 = n280 ;
  assign y191 = n281 ;
  assign y192 = n283 ;
  assign y193 = n284 ;
  assign y194 = n285 ;
  assign y195 = n286 ;
  assign y196 = n287 ;
  assign y197 = n288 ;
  assign y198 = n289 ;
  assign y199 = n290 ;
  assign y200 = n291 ;
  assign y201 = n292 ;
  assign y202 = n293 ;
  assign y203 = n294 ;
  assign y204 = n295 ;
  assign y205 = n296 ;
  assign y206 = n297 ;
  assign y207 = n298 ;
  assign y208 = n300 ;
  assign y209 = n301 ;
  assign y210 = n302 ;
  assign y211 = n303 ;
  assign y212 = n304 ;
  assign y213 = n305 ;
  assign y214 = n306 ;
  assign y215 = n307 ;
  assign y216 = n308 ;
  assign y217 = n309 ;
  assign y218 = n310 ;
  assign y219 = n311 ;
  assign y220 = n312 ;
  assign y221 = n313 ;
  assign y222 = n314 ;
  assign y223 = n315 ;
  assign y224 = n317 ;
  assign y225 = n318 ;
  assign y226 = n319 ;
  assign y227 = n320 ;
  assign y228 = n321 ;
  assign y229 = n322 ;
  assign y230 = n323 ;
  assign y231 = n324 ;
  assign y232 = n325 ;
  assign y233 = n326 ;
  assign y234 = n327 ;
  assign y235 = n328 ;
  assign y236 = n329 ;
  assign y237 = n330 ;
  assign y238 = n331 ;
  assign y239 = n332 ;
  assign y240 = n334 ;
  assign y241 = n335 ;
  assign y242 = n336 ;
  assign y243 = n337 ;
  assign y244 = n338 ;
  assign y245 = n339 ;
  assign y246 = n340 ;
  assign y247 = n341 ;
  assign y248 = n342 ;
  assign y249 = n343 ;
  assign y250 = n344 ;
  assign y251 = n345 ;
  assign y252 = n346 ;
  assign y253 = n347 ;
  assign y254 = n348 ;
  assign y255 = n349 ;
endmodule
