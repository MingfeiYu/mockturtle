module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n802 , n803 , n804 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n823 , n824 , n825 , n826 , n827 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n999 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1164 , n1165 , n1166 , n1169 , n1170 , n1171 , n1172 , n1173 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1216 , n1217 , n1218 , n1221 , n1222 , n1223 , n1224 , n1225 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1268 , n1269 , n1270 , n1273 , n1274 , n1275 , n1276 , n1277 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1422 , n1423 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1593 , n1594 , n1597 , n1598 , n1599 , n1600 , n1601 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1640 , n1641 , n1642 , n1645 , n1646 , n1647 , n1648 , n1649 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1793 , n1794 , n1795 , n1798 , n1799 , n1800 , n1801 , n1802 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1947 , n1948 , n1951 , n1952 , n1953 , n1954 , n1955 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2123 , n2124 , n2127 , n2128 , n2129 , n2130 , n2131 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2262 , n2263 , n2264 , n2265 ;
  assign n257 = ~x129 & ~x130 ;
  assign n258 = x1 & n257 ;
  assign n259 = x2 & ~x3 ;
  assign n260 = ~x130 & n259 ;
  assign n261 = n260 ^ x3 ;
  assign n262 = n258 & ~n261 ;
  assign n263 = n262 ^ n261 ;
  assign n264 = ~x131 & ~x132 ;
  assign n265 = x4 & ~x5 ;
  assign n266 = ~x132 & n265 ;
  assign n267 = n266 ^ x5 ;
  assign n268 = n264 & ~n267 ;
  assign n269 = n263 & n268 ;
  assign n270 = n269 ^ n267 ;
  assign n271 = ~x252 & ~x253 ;
  assign n272 = ~x254 & n271 ;
  assign n273 = ~x221 & ~x222 ;
  assign n274 = ~x248 & ~x250 ;
  assign n275 = ~x249 & n274 ;
  assign n276 = ~x247 & ~x251 ;
  assign n277 = n275 & n276 ;
  assign n278 = ~x246 & n277 ;
  assign n279 = ~x245 & n278 ;
  assign n280 = ~x241 & ~x242 ;
  assign n281 = ~x240 & n280 ;
  assign n282 = ~x243 & n281 ;
  assign n283 = ~x244 & n282 ;
  assign n284 = n279 & n283 ;
  assign n285 = ~x238 & ~x239 ;
  assign n286 = n284 & n285 ;
  assign n287 = ~x235 & ~x237 ;
  assign n288 = ~x236 & n287 ;
  assign n289 = ~x229 & ~x230 ;
  assign n290 = ~x228 & n289 ;
  assign n291 = ~x231 & n290 ;
  assign n292 = ~x227 & ~x232 ;
  assign n293 = n291 & n292 ;
  assign n294 = ~x226 & ~x233 ;
  assign n295 = n293 & n294 ;
  assign n296 = ~x234 & n295 ;
  assign n297 = n288 & n296 ;
  assign n298 = n286 & n297 ;
  assign n299 = ~x224 & ~x225 ;
  assign n300 = ~x223 & n299 ;
  assign n301 = n298 & n300 ;
  assign n302 = n273 & n301 ;
  assign n303 = ~x216 & ~x217 ;
  assign n304 = ~x218 & n303 ;
  assign n305 = ~x219 & n304 ;
  assign n306 = ~x212 & ~x213 ;
  assign n307 = ~x214 & n306 ;
  assign n308 = ~x215 & n307 ;
  assign n309 = ~x209 & ~x210 ;
  assign n310 = ~x208 & n309 ;
  assign n311 = ~x211 & n310 ;
  assign n312 = n308 & n311 ;
  assign n313 = n305 & n312 ;
  assign n314 = ~x205 & ~x206 ;
  assign n315 = ~x207 & n314 ;
  assign n316 = ~x203 & ~x204 ;
  assign n317 = n315 & n316 ;
  assign n318 = ~x200 & ~x202 ;
  assign n319 = ~x201 & n318 ;
  assign n320 = n317 & n319 ;
  assign n321 = n313 & n320 ;
  assign n322 = ~x220 & n321 ;
  assign n323 = n302 & n322 ;
  assign n324 = ~x197 & ~x198 ;
  assign n325 = ~x196 & n324 ;
  assign n326 = ~x199 & n325 ;
  assign n327 = ~x193 & ~x194 ;
  assign n328 = ~x192 & n327 ;
  assign n329 = ~x195 & n328 ;
  assign n330 = n326 & n329 ;
  assign n331 = ~x188 & ~x189 ;
  assign n332 = ~x190 & n331 ;
  assign n333 = ~x191 & n332 ;
  assign n334 = ~x184 & ~x185 ;
  assign n335 = ~x186 & n334 ;
  assign n336 = ~x187 & n335 ;
  assign n337 = n333 & n336 ;
  assign n338 = n330 & n337 ;
  assign n339 = n323 & n338 ;
  assign n340 = ~x180 & ~x181 ;
  assign n341 = ~x182 & n340 ;
  assign n342 = ~x183 & n341 ;
  assign n343 = ~x176 & ~x178 ;
  assign n344 = ~x177 & n343 ;
  assign n345 = ~x179 & n344 ;
  assign n346 = n342 & n345 ;
  assign n347 = n339 & n346 ;
  assign n348 = n272 & n347 ;
  assign n349 = ~x173 & ~x174 ;
  assign n350 = ~x172 & n349 ;
  assign n351 = ~x171 & ~x175 ;
  assign n352 = n350 & n351 ;
  assign n353 = ~x170 & n352 ;
  assign n354 = ~x168 & ~x169 ;
  assign n355 = n353 & n354 ;
  assign n356 = n348 & n355 ;
  assign n357 = ~x165 & ~x166 ;
  assign n358 = ~x164 & n357 ;
  assign n359 = ~x167 & n358 ;
  assign n360 = n356 & n359 ;
  assign n361 = ~x161 & ~x162 ;
  assign n362 = ~x160 & n361 ;
  assign n363 = ~x163 & n362 ;
  assign n364 = n360 & n363 ;
  assign n365 = ~x157 & ~x158 ;
  assign n366 = ~x156 & n365 ;
  assign n367 = ~x159 & n366 ;
  assign n368 = n364 & n367 ;
  assign n369 = ~x154 & ~x155 ;
  assign n370 = n368 & n369 ;
  assign n371 = ~x153 & n370 ;
  assign n372 = ~x150 & ~x151 ;
  assign n373 = ~x149 & n372 ;
  assign n374 = ~x147 & ~x148 ;
  assign n375 = n373 & n374 ;
  assign n376 = ~x146 & ~x152 ;
  assign n377 = n375 & n376 ;
  assign n378 = n371 & n377 ;
  assign n379 = ~x142 & ~x144 ;
  assign n380 = ~x143 & n379 ;
  assign n381 = ~x145 & n380 ;
  assign n382 = ~x141 & n381 ;
  assign n383 = n378 & n382 ;
  assign n384 = ~x139 & ~x140 ;
  assign n385 = ~x138 & n384 ;
  assign n386 = n383 & n385 ;
  assign n387 = ~x134 & ~x135 ;
  assign n388 = ~x136 & n387 ;
  assign n389 = ~x133 & ~x137 ;
  assign n390 = n388 & n389 ;
  assign n391 = ~x255 & n390 ;
  assign n392 = n386 & n391 ;
  assign n393 = x12 & ~x140 ;
  assign n394 = ~x13 & ~n393 ;
  assign n395 = x11 & n384 ;
  assign n396 = n394 & n395 ;
  assign n397 = n396 ^ n394 ;
  assign n398 = x14 & n381 ;
  assign n399 = ~x18 & ~x145 ;
  assign n400 = ~x16 & ~x144 ;
  assign n408 = x15 & n400 ;
  assign n409 = ~x143 & n408 ;
  assign n410 = n409 ^ x143 ;
  assign n401 = n400 ^ x144 ;
  assign n402 = n401 ^ x143 ;
  assign n411 = n410 ^ n402 ;
  assign n412 = ~x17 & n411 ;
  assign n413 = n399 & ~n412 ;
  assign n414 = n413 ^ x18 ;
  assign n415 = n398 & ~n414 ;
  assign n416 = n415 ^ n414 ;
  assign n417 = x26 & n370 ;
  assign n418 = x27 & ~x28 ;
  assign n419 = ~x155 & n418 ;
  assign n420 = n419 ^ x28 ;
  assign n421 = x29 & n365 ;
  assign n422 = x30 & ~x31 ;
  assign n423 = ~x158 & n422 ;
  assign n424 = n423 ^ x31 ;
  assign n425 = n421 & ~n424 ;
  assign n426 = n425 ^ n424 ;
  assign n427 = ~x32 & ~x159 ;
  assign n428 = n426 & n427 ;
  assign n429 = n428 ^ x32 ;
  assign n430 = x33 & n361 ;
  assign n431 = x34 & ~x35 ;
  assign n432 = ~x162 & n431 ;
  assign n433 = n432 ^ x35 ;
  assign n434 = n430 & ~n433 ;
  assign n435 = n434 ^ n433 ;
  assign n436 = ~x36 & ~x163 ;
  assign n437 = n435 & n436 ;
  assign n438 = n437 ^ x36 ;
  assign n439 = x37 & n357 ;
  assign n440 = x38 & ~x39 ;
  assign n441 = ~x166 & n440 ;
  assign n442 = n441 ^ x39 ;
  assign n443 = n439 & ~n442 ;
  assign n444 = n443 ^ n442 ;
  assign n445 = ~x40 & ~x167 ;
  assign n446 = n444 & n445 ;
  assign n447 = n446 ^ x40 ;
  assign n448 = x41 & ~x42 ;
  assign n449 = ~x169 & n448 ;
  assign n450 = n449 ^ x42 ;
  assign n451 = x45 & n349 ;
  assign n452 = x46 & ~x47 ;
  assign n453 = ~x174 & n452 ;
  assign n454 = n453 ^ x47 ;
  assign n455 = n451 & ~n454 ;
  assign n456 = n455 ^ n454 ;
  assign n457 = ~x175 & ~n456 ;
  assign n458 = n350 & n457 ;
  assign n459 = x44 & n458 ;
  assign n460 = n459 ^ n457 ;
  assign n461 = n460 ^ x175 ;
  assign n462 = ~x48 & n461 ;
  assign n463 = x43 & n352 ;
  assign n464 = n462 & n463 ;
  assign n465 = n464 ^ n462 ;
  assign n466 = n353 & n465 ;
  assign n467 = n450 & n466 ;
  assign n468 = n467 ^ n465 ;
  assign n469 = ~x52 & ~x179 ;
  assign n470 = ~x50 & ~x178 ;
  assign n478 = x49 & n470 ;
  assign n479 = ~x177 & n478 ;
  assign n480 = n479 ^ x177 ;
  assign n471 = n470 ^ x178 ;
  assign n472 = n471 ^ x177 ;
  assign n481 = n480 ^ n472 ;
  assign n482 = ~x51 & n481 ;
  assign n483 = n469 & ~n482 ;
  assign n484 = n483 ^ x52 ;
  assign n485 = x53 & ~x54 ;
  assign n486 = ~x181 & n485 ;
  assign n487 = n486 ^ x54 ;
  assign n488 = ~x55 & ~x182 ;
  assign n489 = n487 & n488 ;
  assign n490 = n489 ^ x55 ;
  assign n491 = ~x56 & ~x183 ;
  assign n492 = n490 & n491 ;
  assign n493 = n492 ^ x56 ;
  assign n494 = n342 & ~n493 ;
  assign n495 = n484 & n494 ;
  assign n496 = n495 ^ n493 ;
  assign n497 = x57 & ~x58 ;
  assign n498 = ~x185 & n497 ;
  assign n499 = n498 ^ x58 ;
  assign n500 = ~x59 & ~x186 ;
  assign n501 = n499 & n500 ;
  assign n502 = n501 ^ x59 ;
  assign n503 = ~x60 & ~x187 ;
  assign n504 = n502 & n503 ;
  assign n505 = n504 ^ x60 ;
  assign n506 = x61 & ~x62 ;
  assign n507 = ~x189 & n506 ;
  assign n508 = n507 ^ x62 ;
  assign n509 = ~x63 & ~x190 ;
  assign n510 = n508 & n509 ;
  assign n511 = n510 ^ x63 ;
  assign n512 = ~x64 & ~x191 ;
  assign n513 = n511 & n512 ;
  assign n514 = n513 ^ x64 ;
  assign n515 = n333 & ~n514 ;
  assign n516 = n505 & n515 ;
  assign n517 = n516 ^ n514 ;
  assign n518 = x65 & n327 ;
  assign n519 = x66 & ~x67 ;
  assign n520 = ~x194 & n519 ;
  assign n521 = n520 ^ x67 ;
  assign n522 = n518 & ~n521 ;
  assign n523 = n522 ^ n521 ;
  assign n524 = ~x68 & ~x195 ;
  assign n525 = n523 & n524 ;
  assign n526 = n525 ^ x68 ;
  assign n527 = x69 & n324 ;
  assign n528 = x70 & ~x71 ;
  assign n529 = ~x198 & n528 ;
  assign n530 = n529 ^ x71 ;
  assign n531 = n527 & ~n530 ;
  assign n532 = n531 ^ n530 ;
  assign n533 = ~x72 & ~x199 ;
  assign n534 = n532 & n533 ;
  assign n535 = n534 ^ x72 ;
  assign n536 = n326 & ~n535 ;
  assign n537 = n526 & n536 ;
  assign n538 = n537 ^ n535 ;
  assign n539 = n330 & ~n538 ;
  assign n540 = n517 & n539 ;
  assign n541 = n540 ^ n538 ;
  assign n542 = x76 & ~x77 ;
  assign n543 = ~x204 & n542 ;
  assign n544 = n543 ^ x77 ;
  assign n545 = x78 & ~x79 ;
  assign n546 = ~x206 & n545 ;
  assign n547 = n546 ^ x79 ;
  assign n548 = ~x80 & ~x207 ;
  assign n549 = n547 & n548 ;
  assign n550 = n549 ^ x80 ;
  assign n551 = n315 & ~n550 ;
  assign n552 = n544 & n551 ;
  assign n553 = n552 ^ n550 ;
  assign n554 = n317 & ~n553 ;
  assign n555 = ~x74 & ~x202 ;
  assign n563 = x73 & n555 ;
  assign n564 = ~x201 & n563 ;
  assign n565 = n564 ^ x201 ;
  assign n556 = n555 ^ x202 ;
  assign n557 = n556 ^ x201 ;
  assign n566 = n565 ^ n557 ;
  assign n567 = ~x75 & n566 ;
  assign n568 = n554 & ~n567 ;
  assign n569 = n568 ^ n553 ;
  assign n570 = x81 & n309 ;
  assign n571 = x82 & ~x83 ;
  assign n572 = ~x210 & n571 ;
  assign n573 = n572 ^ x83 ;
  assign n574 = n570 & ~n573 ;
  assign n575 = n574 ^ n573 ;
  assign n576 = ~x84 & ~x211 ;
  assign n577 = n575 & n576 ;
  assign n578 = n577 ^ x84 ;
  assign n579 = x85 & ~x86 ;
  assign n580 = ~x213 & n579 ;
  assign n581 = n580 ^ x86 ;
  assign n582 = ~x87 & ~x214 ;
  assign n583 = n581 & n582 ;
  assign n584 = n583 ^ x87 ;
  assign n585 = ~x88 & ~x215 ;
  assign n586 = n584 & n585 ;
  assign n587 = n586 ^ x88 ;
  assign n588 = n308 & ~n587 ;
  assign n589 = n578 & n588 ;
  assign n590 = n589 ^ n587 ;
  assign n591 = x89 & ~x90 ;
  assign n592 = ~x217 & n591 ;
  assign n593 = n592 ^ x90 ;
  assign n594 = ~x91 & ~x218 ;
  assign n595 = n593 & n594 ;
  assign n596 = n595 ^ x91 ;
  assign n597 = ~x92 & ~x219 ;
  assign n598 = n596 & n597 ;
  assign n599 = n598 ^ x92 ;
  assign n600 = n305 & ~n599 ;
  assign n601 = n590 & n600 ;
  assign n602 = n601 ^ n599 ;
  assign n603 = n313 & ~n602 ;
  assign n604 = n569 & n603 ;
  assign n605 = n604 ^ n602 ;
  assign n606 = ~x220 & n605 ;
  assign n607 = n302 & n606 ;
  assign n608 = x96 & n299 ;
  assign n609 = x97 & ~x98 ;
  assign n610 = ~x225 & n609 ;
  assign n611 = n610 ^ x98 ;
  assign n612 = n608 & ~n611 ;
  assign n613 = n612 ^ n611 ;
  assign n614 = ~n300 & ~n613 ;
  assign n615 = n298 & ~n614 ;
  assign n616 = ~x109 & ~x237 ;
  assign n617 = ~x236 & n616 ;
  assign n618 = x108 & n617 ;
  assign n619 = n618 ^ n616 ;
  assign n620 = n619 ^ x237 ;
  assign n621 = ~x110 & n620 ;
  assign n622 = ~x107 & ~x234 ;
  assign n623 = x101 & n289 ;
  assign n624 = x102 & ~x103 ;
  assign n625 = ~x230 & n624 ;
  assign n626 = n625 ^ x103 ;
  assign n627 = n623 & ~n626 ;
  assign n628 = n627 ^ n626 ;
  assign n629 = ~x104 & ~x231 ;
  assign n630 = n628 & n629 ;
  assign n631 = n630 ^ x104 ;
  assign n632 = ~x232 & ~n631 ;
  assign n640 = n291 & n632 ;
  assign n641 = x100 & n640 ;
  assign n642 = n641 ^ x100 ;
  assign n633 = n632 ^ x232 ;
  assign n634 = n633 ^ x100 ;
  assign n643 = n642 ^ n634 ;
  assign n644 = ~x105 & n643 ;
  assign n645 = ~x233 & n644 ;
  assign n653 = n293 & n645 ;
  assign n654 = x99 & n653 ;
  assign n655 = n654 ^ x99 ;
  assign n646 = n645 ^ x233 ;
  assign n647 = n646 ^ x99 ;
  assign n656 = n655 ^ n647 ;
  assign n657 = ~x106 & n656 ;
  assign n658 = n622 & ~n657 ;
  assign n659 = n658 ^ x107 ;
  assign n660 = n288 & n659 ;
  assign n661 = n621 & n660 ;
  assign n662 = n661 ^ n621 ;
  assign n663 = x111 & ~x112 ;
  assign n664 = ~x239 & n663 ;
  assign n665 = n664 ^ x112 ;
  assign n666 = x113 & n280 ;
  assign n667 = x114 & ~x115 ;
  assign n668 = ~x242 & n667 ;
  assign n669 = n668 ^ x115 ;
  assign n670 = n666 & ~n669 ;
  assign n671 = n670 ^ n669 ;
  assign n672 = ~x116 & ~x243 ;
  assign n673 = n671 & n672 ;
  assign n674 = n673 ^ x116 ;
  assign n675 = ~x117 & ~x244 ;
  assign n676 = n674 & n675 ;
  assign n677 = n676 ^ x117 ;
  assign n678 = x118 & n278 ;
  assign n679 = ~x122 & ~x250 ;
  assign n687 = x121 & n679 ;
  assign n688 = ~x249 & n687 ;
  assign n689 = n688 ^ x249 ;
  assign n680 = n679 ^ x250 ;
  assign n681 = n680 ^ x249 ;
  assign n690 = n689 ^ n681 ;
  assign n691 = ~x123 & n690 ;
  assign n692 = ~x251 & n691 ;
  assign n700 = n275 & n692 ;
  assign n701 = x120 & n700 ;
  assign n702 = n701 ^ x120 ;
  assign n693 = n692 ^ x251 ;
  assign n694 = n693 ^ x120 ;
  assign n703 = n702 ^ n694 ;
  assign n704 = ~x124 & n703 ;
  assign n705 = x119 & n277 ;
  assign n706 = n704 & n705 ;
  assign n707 = n706 ^ n704 ;
  assign n708 = n678 & n707 ;
  assign n709 = n708 ^ n707 ;
  assign n710 = n279 & n709 ;
  assign n711 = n677 & n710 ;
  assign n712 = n711 ^ n709 ;
  assign n713 = n284 & n712 ;
  assign n714 = n665 & n713 ;
  assign n715 = n714 ^ n712 ;
  assign n716 = n286 & n715 ;
  assign n717 = ~n662 & n716 ;
  assign n718 = n717 ^ n715 ;
  assign n719 = ~x96 & ~x97 ;
  assign n720 = x94 & ~x222 ;
  assign n721 = ~x95 & ~n720 ;
  assign n722 = ~x98 & n721 ;
  assign n723 = n719 & n722 ;
  assign n724 = x93 & n273 ;
  assign n725 = n723 & n724 ;
  assign n726 = n725 ^ n723 ;
  assign n727 = n718 & ~n726 ;
  assign n728 = n615 & n727 ;
  assign n729 = n728 ^ n718 ;
  assign n730 = n607 & n729 ;
  assign n731 = n730 ^ n729 ;
  assign n732 = n323 & n731 ;
  assign n733 = n541 & n732 ;
  assign n734 = n733 ^ n731 ;
  assign n735 = n339 & n734 ;
  assign n736 = n496 & n735 ;
  assign n737 = n736 ^ n734 ;
  assign n738 = x125 & ~x126 ;
  assign n739 = ~x253 & n738 ;
  assign n740 = n739 ^ x126 ;
  assign n741 = ~x127 & ~x254 ;
  assign n742 = n740 & n741 ;
  assign n743 = n742 ^ x127 ;
  assign n744 = n272 & ~n743 ;
  assign n745 = ~n737 & n744 ;
  assign n746 = n745 ^ n743 ;
  assign n747 = n348 & ~n746 ;
  assign n748 = ~n468 & n747 ;
  assign n749 = n748 ^ n746 ;
  assign n750 = n356 & ~n749 ;
  assign n751 = n447 & n750 ;
  assign n752 = n751 ^ n749 ;
  assign n753 = n360 & ~n752 ;
  assign n754 = n438 & n753 ;
  assign n755 = n754 ^ n752 ;
  assign n756 = n364 & ~n755 ;
  assign n757 = n429 & n756 ;
  assign n758 = n757 ^ n755 ;
  assign n759 = n368 & ~n758 ;
  assign n760 = n420 & n759 ;
  assign n761 = n760 ^ n758 ;
  assign n762 = n417 & ~n761 ;
  assign n763 = n762 ^ n761 ;
  assign n764 = n371 & ~n763 ;
  assign n765 = x20 & ~x148 ;
  assign n766 = n373 & n765 ;
  assign n767 = x21 & n373 ;
  assign n768 = x22 & n372 ;
  assign n769 = x23 & ~x24 ;
  assign n770 = ~x151 & n769 ;
  assign n771 = n770 ^ x24 ;
  assign n772 = n768 & ~n771 ;
  assign n773 = n772 ^ n771 ;
  assign n774 = n767 & ~n773 ;
  assign n775 = n774 ^ n773 ;
  assign n776 = ~x152 & ~n775 ;
  assign n777 = ~n766 & n776 ;
  assign n785 = n375 & n777 ;
  assign n786 = x19 & n785 ;
  assign n787 = n786 ^ x19 ;
  assign n778 = n777 ^ x152 ;
  assign n779 = n778 ^ x19 ;
  assign n788 = n787 ^ n779 ;
  assign n789 = ~x25 & n788 ;
  assign n790 = n764 & ~n789 ;
  assign n791 = n790 ^ n763 ;
  assign n792 = n378 & ~n791 ;
  assign n793 = n416 & n792 ;
  assign n794 = n793 ^ n791 ;
  assign n795 = n383 & ~n794 ;
  assign n796 = ~n397 & n795 ;
  assign n797 = n796 ^ n794 ;
  assign n798 = ~x255 & ~n797 ;
  assign n802 = ~x8 & ~x136 ;
  assign n810 = x7 & n802 ;
  assign n811 = ~x135 & n810 ;
  assign n812 = n811 ^ x135 ;
  assign n803 = n802 ^ x136 ;
  assign n804 = n803 ^ x135 ;
  assign n813 = n812 ^ n804 ;
  assign n814 = ~x9 & n813 ;
  assign n815 = ~x137 & n814 ;
  assign n823 = n388 & n815 ;
  assign n824 = x6 & n823 ;
  assign n825 = n824 ^ x6 ;
  assign n816 = n815 ^ x137 ;
  assign n817 = n816 ^ x6 ;
  assign n826 = n825 ^ n817 ;
  assign n827 = ~x10 & n826 ;
  assign n832 = n798 & ~n827 ;
  assign n833 = n386 & n832 ;
  assign n834 = n833 ^ n386 ;
  assign n799 = n798 ^ x255 ;
  assign n800 = n799 ^ n386 ;
  assign n835 = n834 ^ n800 ;
  assign n836 = ~x0 & n835 ;
  assign n837 = x128 & n836 ;
  assign n838 = n392 & n837 ;
  assign n839 = n270 & n838 ;
  assign n840 = n839 ^ n837 ;
  assign n841 = n840 ^ x128 ;
  assign n842 = n392 & n836 ;
  assign n847 = n261 & n268 ;
  assign n848 = n847 ^ n267 ;
  assign n849 = n842 & n848 ;
  assign n850 = n849 ^ n836 ;
  assign n851 = ~x128 & ~n850 ;
  assign n852 = ~x1 & ~n851 ;
  assign n853 = x129 & ~n852 ;
  assign n854 = ~n267 & n392 ;
  assign n862 = x3 & n854 ;
  assign n863 = n264 & n862 ;
  assign n864 = n863 ^ n264 ;
  assign n855 = n854 ^ n392 ;
  assign n856 = n855 ^ n264 ;
  assign n865 = n864 ^ n856 ;
  assign n866 = n836 & ~n865 ;
  assign n867 = ~x128 & ~n866 ;
  assign n868 = ~x1 & ~n867 ;
  assign n869 = ~x2 & x130 ;
  assign n870 = ~x129 & n869 ;
  assign n871 = ~n868 & n870 ;
  assign n872 = n871 ^ n869 ;
  assign n873 = n872 ^ x130 ;
  assign n874 = ~x128 & n257 ;
  assign n875 = x131 & ~n263 ;
  assign n876 = ~n868 & n875 ;
  assign n877 = n874 & n876 ;
  assign n878 = n877 ^ n875 ;
  assign n879 = n878 ^ x131 ;
  assign n880 = n836 & n874 ;
  assign n888 = x5 & n880 ;
  assign n889 = n392 & n888 ;
  assign n890 = n889 ^ n392 ;
  assign n881 = n880 ^ n874 ;
  assign n882 = n881 ^ n392 ;
  assign n891 = n890 ^ n882 ;
  assign n892 = ~n263 & ~n891 ;
  assign n893 = ~x131 & ~n892 ;
  assign n894 = ~x4 & ~n893 ;
  assign n895 = x132 & ~n894 ;
  assign n896 = n264 & n874 ;
  assign n897 = ~n270 & n896 ;
  assign n898 = ~n836 & n897 ;
  assign n899 = n898 ^ n270 ;
  assign n900 = ~x133 & n899 ;
  assign n901 = n900 ^ n899 ;
  assign n902 = ~x6 & ~n900 ;
  assign n903 = ~x134 & ~n902 ;
  assign n904 = n903 ^ n902 ;
  assign n905 = ~x7 & ~n903 ;
  assign n906 = ~x135 & ~n905 ;
  assign n907 = n906 ^ n905 ;
  assign n908 = ~x8 & x136 ;
  assign n909 = ~n906 & n908 ;
  assign n910 = n909 ^ x136 ;
  assign n911 = x137 & n814 ;
  assign n912 = ~n902 & n911 ;
  assign n913 = n388 & n912 ;
  assign n914 = n913 ^ n911 ;
  assign n915 = n914 ^ x137 ;
  assign n916 = n391 & n896 ;
  assign n917 = ~n270 & n390 ;
  assign n925 = x0 & n917 ;
  assign n926 = n896 & n925 ;
  assign n927 = n926 ^ n896 ;
  assign n918 = n917 ^ n390 ;
  assign n919 = n918 ^ n896 ;
  assign n928 = n927 ^ n919 ;
  assign n929 = n827 & ~n928 ;
  assign n930 = x138 & n929 ;
  assign n931 = n916 & n930 ;
  assign n932 = n797 & n931 ;
  assign n933 = n932 ^ n930 ;
  assign n934 = n933 ^ x138 ;
  assign n935 = ~x138 & n916 ;
  assign n936 = ~n794 & n935 ;
  assign n944 = x13 & n936 ;
  assign n945 = n383 & n944 ;
  assign n946 = n945 ^ n383 ;
  assign n937 = n936 ^ n935 ;
  assign n938 = n937 ^ n383 ;
  assign n947 = n946 ^ n938 ;
  assign n948 = ~x11 & ~n947 ;
  assign n949 = ~x138 & ~n929 ;
  assign n950 = n948 & n949 ;
  assign n951 = n950 ^ n948 ;
  assign n952 = n393 & n935 ;
  assign n953 = n383 & n952 ;
  assign n954 = n953 ^ x139 ;
  assign n955 = x139 & n954 ;
  assign n956 = n951 & n955 ;
  assign n957 = n956 ^ x139 ;
  assign n958 = ~x12 & x140 ;
  assign n959 = ~x139 & n958 ;
  assign n960 = ~n951 & n959 ;
  assign n961 = n960 ^ n958 ;
  assign n962 = n961 ^ x140 ;
  assign n963 = n385 & n916 ;
  assign n964 = n385 & n397 ;
  assign n965 = ~n929 & n964 ;
  assign n966 = n965 ^ n397 ;
  assign n967 = x141 & n966 ;
  assign n968 = n963 & n967 ;
  assign n969 = n794 & n968 ;
  assign n970 = n969 ^ n967 ;
  assign n971 = n970 ^ x141 ;
  assign n972 = ~x141 & n378 ;
  assign n973 = n963 & n972 ;
  assign n974 = n963 ^ x141 ;
  assign n975 = n974 ^ x14 ;
  assign n976 = n966 ^ n963 ;
  assign n977 = n976 ^ x14 ;
  assign n978 = n966 ^ n791 ;
  assign n979 = n978 ^ x141 ;
  assign n980 = ~n977 & ~n979 ;
  assign n981 = n975 & n980 ;
  assign n982 = n981 ^ n966 ;
  assign n983 = n982 ^ x141 ;
  assign n984 = ~x14 & ~n983 ;
  assign n985 = ~x141 & n984 ;
  assign n986 = n985 ^ x14 ;
  assign n987 = x142 & ~n986 ;
  assign n988 = n973 & n987 ;
  assign n989 = n414 & n988 ;
  assign n990 = n989 ^ n987 ;
  assign n991 = n990 ^ x142 ;
  assign n992 = x18 & n973 ;
  assign n993 = ~n986 & n992 ;
  assign n994 = n993 ^ n986 ;
  assign n995 = ~x142 & ~n994 ;
  assign n999 = ~x145 & n973 ;
  assign n1004 = n995 & n999 ;
  assign n1005 = x17 & n1004 ;
  assign n1006 = n1005 ^ x17 ;
  assign n996 = n995 ^ x142 ;
  assign n997 = n996 ^ x17 ;
  assign n1007 = n1006 ^ n997 ;
  assign n1008 = ~x15 & n1007 ;
  assign n1009 = n379 & n999 ;
  assign n1010 = x16 & n1009 ;
  assign n1011 = n1010 ^ x143 ;
  assign n1012 = x143 & n1011 ;
  assign n1013 = n1008 & n1012 ;
  assign n1014 = n1013 ^ x143 ;
  assign n1015 = ~x16 & x144 ;
  assign n1016 = ~x143 & n1015 ;
  assign n1017 = ~n1008 & n1016 ;
  assign n1018 = n1017 ^ n1015 ;
  assign n1019 = n1018 ^ x144 ;
  assign n1020 = x145 & n412 ;
  assign n1021 = n994 & n1020 ;
  assign n1022 = n380 & n1021 ;
  assign n1023 = n1022 ^ n1020 ;
  assign n1024 = n1023 ^ x145 ;
  assign n1025 = x146 & ~n414 ;
  assign n1026 = n381 & n1025 ;
  assign n1027 = n986 & n1026 ;
  assign n1028 = n1027 ^ n1025 ;
  assign n1029 = n1028 ^ x146 ;
  assign n1030 = n382 & n963 ;
  assign n1031 = n371 & n376 ;
  assign n1032 = n1030 & n1031 ;
  assign n1033 = n382 & ~n416 ;
  assign n1034 = ~n966 & n1033 ;
  assign n1035 = n1034 ^ n416 ;
  assign n1036 = ~n763 & n1030 ;
  assign n1044 = x25 & n1036 ;
  assign n1045 = n371 & n1044 ;
  assign n1046 = n1045 ^ n371 ;
  assign n1037 = n1036 ^ n1030 ;
  assign n1038 = n1037 ^ n371 ;
  assign n1047 = n1046 ^ n1038 ;
  assign n1048 = ~n1035 & ~n1047 ;
  assign n1049 = ~x146 & ~n1048 ;
  assign n1050 = ~x19 & ~n1049 ;
  assign n1051 = n775 & n1032 ;
  assign n1052 = n1050 & n1051 ;
  assign n1053 = n1052 ^ n1050 ;
  assign n1054 = x147 & n1053 ;
  assign n1055 = n1032 & n1054 ;
  assign n1056 = n766 & n1055 ;
  assign n1057 = n1056 ^ n1054 ;
  assign n1058 = n1057 ^ x147 ;
  assign n1059 = ~x20 & x148 ;
  assign n1060 = ~x147 & n1059 ;
  assign n1061 = ~n1053 & n1060 ;
  assign n1062 = n1061 ^ n1059 ;
  assign n1063 = n1062 ^ x148 ;
  assign n1064 = n374 & n1032 ;
  assign n1065 = ~x21 & ~n765 ;
  assign n1066 = n374 & ~n1050 ;
  assign n1067 = n1065 & n1066 ;
  assign n1068 = n1067 ^ n1065 ;
  assign n1069 = x149 & n1068 ;
  assign n1070 = n1064 & n1069 ;
  assign n1071 = n773 & n1070 ;
  assign n1072 = n1071 ^ n1069 ;
  assign n1073 = n1072 ^ x149 ;
  assign n1074 = ~x149 & n1068 ;
  assign n1082 = n771 & n1074 ;
  assign n1083 = n1064 & n1082 ;
  assign n1084 = n1083 ^ n1064 ;
  assign n1075 = n1074 ^ x149 ;
  assign n1076 = n1075 ^ n1064 ;
  assign n1085 = n1084 ^ n1076 ;
  assign n1086 = ~x22 & n1085 ;
  assign n1087 = x150 & ~n1086 ;
  assign n1090 = n1064 & n1074 ;
  assign n1091 = x24 & n1090 ;
  assign n1092 = n1091 ^ x24 ;
  assign n1088 = n1075 ^ x24 ;
  assign n1093 = n1092 ^ n1088 ;
  assign n1094 = ~x22 & n1093 ;
  assign n1095 = ~x150 & ~n1094 ;
  assign n1096 = ~x23 & ~n1095 ;
  assign n1097 = x151 & ~n1096 ;
  assign n1098 = x152 & ~n773 ;
  assign n1099 = n373 & n1098 ;
  assign n1100 = ~n1068 & n1099 ;
  assign n1101 = n1100 ^ n1098 ;
  assign n1102 = n1101 ^ x152 ;
  assign n1103 = n377 & n1030 ;
  assign n1104 = n377 & n1035 ;
  assign n1105 = n789 & n1104 ;
  assign n1106 = n1105 ^ n789 ;
  assign n1107 = x153 & n1106 ;
  assign n1108 = n1103 & n1107 ;
  assign n1109 = n763 & n1108 ;
  assign n1110 = n1109 ^ n1107 ;
  assign n1111 = n1110 ^ x153 ;
  assign n1112 = ~x153 & n1103 ;
  assign n1113 = ~x26 & ~x153 ;
  assign n1114 = ~n1106 & n1113 ;
  assign n1115 = n1114 ^ x26 ;
  assign n1116 = x154 & ~n1115 ;
  assign n1117 = n1112 & n1116 ;
  assign n1118 = n761 & n1117 ;
  assign n1119 = n1118 ^ n1116 ;
  assign n1120 = n1119 ^ x154 ;
  assign n1121 = ~n758 & n1112 ;
  assign n1129 = x28 & n1121 ;
  assign n1130 = n368 & n1129 ;
  assign n1131 = n1130 ^ n368 ;
  assign n1122 = n1121 ^ n1112 ;
  assign n1123 = n1122 ^ n368 ;
  assign n1132 = n1131 ^ n1123 ;
  assign n1133 = ~n1115 & ~n1132 ;
  assign n1134 = ~x154 & ~n1133 ;
  assign n1135 = ~x27 & ~n1134 ;
  assign n1136 = x155 & ~n1135 ;
  assign n1137 = n369 & n1112 ;
  assign n1138 = n369 & ~n420 ;
  assign n1139 = n1115 & n1138 ;
  assign n1140 = n1139 ^ n420 ;
  assign n1141 = x156 & ~n1140 ;
  assign n1142 = n1137 & n1141 ;
  assign n1143 = n758 & n1142 ;
  assign n1144 = n1143 ^ n1141 ;
  assign n1145 = n1144 ^ x156 ;
  assign n1146 = ~x29 & x157 ;
  assign n1164 = ~x159 & n364 ;
  assign n1147 = ~n755 & n1137 ;
  assign n1155 = x32 & n1147 ;
  assign n1156 = n364 & n1155 ;
  assign n1157 = n1156 ^ n364 ;
  assign n1148 = n1147 ^ n1137 ;
  assign n1149 = n1148 ^ n364 ;
  assign n1158 = n1157 ^ n1149 ;
  assign n1159 = ~n1140 & ~n1158 ;
  assign n1160 = ~x156 & n1159 ;
  assign n1165 = n1137 & n1160 ;
  assign n1166 = n1164 & n1165 ;
  assign n1169 = n424 & n1166 ;
  assign n1161 = n1160 ^ x156 ;
  assign n1170 = n1169 ^ n1161 ;
  assign n1171 = n1146 & n1170 ;
  assign n1172 = n1171 ^ x157 ;
  assign n1173 = ~x29 & ~x157 ;
  assign n1178 = x31 & n1166 ;
  assign n1179 = n1178 ^ n1161 ;
  assign n1180 = n1173 & n1179 ;
  assign n1181 = n1180 ^ x157 ;
  assign n1182 = ~x30 & n1181 ;
  assign n1183 = x158 & ~n1182 ;
  assign n1184 = x159 & ~n426 ;
  assign n1185 = n366 & n1184 ;
  assign n1186 = ~n1159 & n1185 ;
  assign n1187 = n1186 ^ n1184 ;
  assign n1188 = n1187 ^ x159 ;
  assign n1189 = n367 & n1137 ;
  assign n1190 = n367 & ~n429 ;
  assign n1191 = n1140 & n1190 ;
  assign n1192 = n1191 ^ n429 ;
  assign n1193 = x160 & ~n1192 ;
  assign n1194 = n1189 & n1193 ;
  assign n1195 = n755 & n1194 ;
  assign n1196 = n1195 ^ n1193 ;
  assign n1197 = n1196 ^ x160 ;
  assign n1198 = ~x33 & x161 ;
  assign n1216 = ~x163 & n360 ;
  assign n1199 = ~n752 & n1189 ;
  assign n1207 = x36 & n1199 ;
  assign n1208 = n360 & n1207 ;
  assign n1209 = n1208 ^ n360 ;
  assign n1200 = n1199 ^ n1189 ;
  assign n1201 = n1200 ^ n360 ;
  assign n1210 = n1209 ^ n1201 ;
  assign n1211 = ~n1192 & ~n1210 ;
  assign n1212 = ~x160 & n1211 ;
  assign n1217 = n1189 & n1212 ;
  assign n1218 = n1216 & n1217 ;
  assign n1221 = n433 & n1218 ;
  assign n1213 = n1212 ^ x160 ;
  assign n1222 = n1221 ^ n1213 ;
  assign n1223 = n1198 & n1222 ;
  assign n1224 = n1223 ^ x161 ;
  assign n1225 = ~x33 & ~x161 ;
  assign n1230 = x35 & n1218 ;
  assign n1231 = n1230 ^ n1213 ;
  assign n1232 = n1225 & n1231 ;
  assign n1233 = n1232 ^ x161 ;
  assign n1234 = ~x34 & n1233 ;
  assign n1235 = x162 & ~n1234 ;
  assign n1236 = x163 & ~n435 ;
  assign n1237 = n362 & n1236 ;
  assign n1238 = ~n1211 & n1237 ;
  assign n1239 = n1238 ^ n1236 ;
  assign n1240 = n1239 ^ x163 ;
  assign n1241 = n363 & n1189 ;
  assign n1242 = n363 & ~n438 ;
  assign n1243 = n1192 & n1242 ;
  assign n1244 = n1243 ^ n438 ;
  assign n1245 = x164 & ~n1244 ;
  assign n1246 = n1241 & n1245 ;
  assign n1247 = n752 & n1246 ;
  assign n1248 = n1247 ^ n1245 ;
  assign n1249 = n1248 ^ x164 ;
  assign n1250 = ~x37 & x165 ;
  assign n1268 = ~x167 & n356 ;
  assign n1251 = ~n749 & n1241 ;
  assign n1259 = x40 & n1251 ;
  assign n1260 = n356 & n1259 ;
  assign n1261 = n1260 ^ n356 ;
  assign n1252 = n1251 ^ n1241 ;
  assign n1253 = n1252 ^ n356 ;
  assign n1262 = n1261 ^ n1253 ;
  assign n1263 = ~n1244 & ~n1262 ;
  assign n1264 = ~x164 & n1263 ;
  assign n1269 = n1241 & n1264 ;
  assign n1270 = n1268 & n1269 ;
  assign n1273 = n442 & n1270 ;
  assign n1265 = n1264 ^ x164 ;
  assign n1274 = n1273 ^ n1265 ;
  assign n1275 = n1250 & n1274 ;
  assign n1276 = n1275 ^ x165 ;
  assign n1277 = ~x37 & ~x165 ;
  assign n1282 = x39 & n1270 ;
  assign n1283 = n1282 ^ n1265 ;
  assign n1284 = n1277 & n1283 ;
  assign n1285 = n1284 ^ x165 ;
  assign n1286 = ~x38 & n1285 ;
  assign n1287 = x166 & ~n1286 ;
  assign n1288 = x167 & ~n444 ;
  assign n1289 = n358 & n1288 ;
  assign n1290 = ~n1263 & n1289 ;
  assign n1291 = n1290 ^ n1288 ;
  assign n1292 = n1291 ^ x167 ;
  assign n1293 = n359 & n1241 ;
  assign n1294 = n359 & ~n447 ;
  assign n1295 = n1244 & n1294 ;
  assign n1296 = n1295 ^ n447 ;
  assign n1297 = x168 & ~n1296 ;
  assign n1298 = n1293 & n1297 ;
  assign n1299 = n749 & n1298 ;
  assign n1300 = n1299 ^ n1297 ;
  assign n1301 = n1300 ^ x168 ;
  assign n1302 = n746 & n1293 ;
  assign n1303 = ~n1296 & n1302 ;
  assign n1304 = n1303 ^ n1296 ;
  assign n1305 = n348 & n1293 ;
  assign n1306 = n465 & n1305 ;
  assign n1314 = n353 & n1306 ;
  assign n1315 = x42 & n1314 ;
  assign n1316 = n1315 ^ x42 ;
  assign n1307 = n1306 ^ n1305 ;
  assign n1308 = n1307 ^ x42 ;
  assign n1317 = n1316 ^ n1308 ;
  assign n1318 = ~n1304 & ~n1317 ;
  assign n1319 = ~x168 & ~n1318 ;
  assign n1320 = ~x41 & ~n1319 ;
  assign n1321 = x169 & ~n1320 ;
  assign n1322 = n354 & n1305 ;
  assign n1323 = n354 & ~n450 ;
  assign n1324 = n1304 & n1323 ;
  assign n1325 = n1324 ^ n450 ;
  assign n1326 = x170 & ~n1325 ;
  assign n1327 = n1322 & n1326 ;
  assign n1328 = ~n465 & n1327 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1330 = n1329 ^ x170 ;
  assign n1331 = ~x170 & n1322 ;
  assign n1332 = n1322 ^ x170 ;
  assign n1333 = n1332 ^ x43 ;
  assign n1334 = n1325 ^ n1322 ;
  assign n1335 = n1334 ^ x43 ;
  assign n1336 = n1325 ^ x48 ;
  assign n1337 = n1336 ^ x170 ;
  assign n1338 = n1335 & n1337 ;
  assign n1339 = n1333 & n1338 ;
  assign n1340 = n1339 ^ n1325 ;
  assign n1341 = n1340 ^ x170 ;
  assign n1342 = ~x43 & n1341 ;
  assign n1343 = ~x170 & n1342 ;
  assign n1344 = n1343 ^ x43 ;
  assign n1345 = x171 & ~n1344 ;
  assign n1346 = n1331 & n1345 ;
  assign n1347 = ~n461 & n1346 ;
  assign n1348 = n1347 ^ n1345 ;
  assign n1349 = n1348 ^ x171 ;
  assign n1350 = n351 & n1331 ;
  assign n1351 = ~x44 & ~x171 ;
  assign n1352 = n1344 & n1351 ;
  assign n1353 = n1352 ^ x44 ;
  assign n1354 = x172 & ~n1353 ;
  assign n1355 = n1350 & n1354 ;
  assign n1356 = n456 & n1355 ;
  assign n1357 = n1356 ^ n1354 ;
  assign n1358 = n1357 ^ x172 ;
  assign n1359 = ~x172 & ~n1353 ;
  assign n1367 = n454 & n1359 ;
  assign n1368 = n1350 & n1367 ;
  assign n1369 = n1368 ^ n1350 ;
  assign n1360 = n1359 ^ x172 ;
  assign n1361 = n1360 ^ n1350 ;
  assign n1370 = n1369 ^ n1361 ;
  assign n1371 = ~x45 & n1370 ;
  assign n1372 = x173 & ~n1371 ;
  assign n1375 = n1350 & n1359 ;
  assign n1376 = x47 & n1375 ;
  assign n1377 = n1376 ^ x47 ;
  assign n1373 = n1360 ^ x47 ;
  assign n1378 = n1377 ^ n1373 ;
  assign n1379 = ~x45 & n1378 ;
  assign n1380 = ~x173 & ~n1379 ;
  assign n1381 = ~x46 & ~n1380 ;
  assign n1382 = x174 & ~n1381 ;
  assign n1383 = x175 & ~n456 ;
  assign n1384 = n350 & n1383 ;
  assign n1385 = n1353 & n1384 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1387 = n1386 ^ x175 ;
  assign n1388 = x176 & n468 ;
  assign n1389 = n355 & n1388 ;
  assign n1390 = n1304 & n1389 ;
  assign n1391 = n1390 ^ n1388 ;
  assign n1392 = n1391 ^ x176 ;
  assign n1393 = n355 & n1293 ;
  assign n1394 = n272 & n1393 ;
  assign n1395 = ~n734 & n1394 ;
  assign n1396 = n743 & n1393 ;
  assign n1397 = n355 & n468 ;
  assign n1398 = n1296 & n1397 ;
  assign n1399 = n1398 ^ n468 ;
  assign n1400 = n1396 & n1399 ;
  assign n1401 = n1400 ^ n1399 ;
  assign n1402 = n1395 & n1401 ;
  assign n1403 = n1402 ^ n1401 ;
  assign n1404 = n339 & n1394 ;
  assign n1405 = ~n493 & n1404 ;
  assign n1413 = n342 & n1405 ;
  assign n1414 = x52 & n1413 ;
  assign n1415 = n1414 ^ x52 ;
  assign n1406 = n1405 ^ n1404 ;
  assign n1407 = n1406 ^ x52 ;
  assign n1416 = n1415 ^ n1407 ;
  assign n1417 = n1403 & ~n1416 ;
  assign n1418 = ~x176 & n1417 ;
  assign n1422 = ~x179 & n342 ;
  assign n1423 = n1404 & n1422 ;
  assign n1428 = n1418 & n1423 ;
  assign n1429 = x51 & n1428 ;
  assign n1430 = n1429 ^ x51 ;
  assign n1419 = n1418 ^ x176 ;
  assign n1420 = n1419 ^ x51 ;
  assign n1431 = n1430 ^ n1420 ;
  assign n1432 = ~x49 & n1431 ;
  assign n1433 = n343 & n1423 ;
  assign n1434 = x50 & n1433 ;
  assign n1435 = n1434 ^ x177 ;
  assign n1436 = x177 & n1435 ;
  assign n1437 = n1432 & n1436 ;
  assign n1438 = n1437 ^ x177 ;
  assign n1439 = ~x50 & x178 ;
  assign n1440 = ~x177 & n1439 ;
  assign n1441 = ~n1432 & n1440 ;
  assign n1442 = n1441 ^ n1439 ;
  assign n1443 = n1442 ^ x178 ;
  assign n1444 = x179 & n482 ;
  assign n1445 = n344 & n1444 ;
  assign n1446 = ~n1417 & n1445 ;
  assign n1447 = n1446 ^ n1444 ;
  assign n1448 = n1447 ^ x179 ;
  assign n1449 = n345 & n1404 ;
  assign n1450 = n345 & ~n484 ;
  assign n1451 = ~n1403 & n1450 ;
  assign n1452 = n1451 ^ n484 ;
  assign n1453 = x180 & ~n1452 ;
  assign n1454 = n1449 & n1453 ;
  assign n1455 = n493 & n1454 ;
  assign n1456 = n1455 ^ n1453 ;
  assign n1457 = n1456 ^ x180 ;
  assign n1458 = ~x183 & n1449 ;
  assign n1459 = x55 & n1458 ;
  assign n1460 = x56 & n1449 ;
  assign n1461 = ~n1452 & n1460 ;
  assign n1462 = n1461 ^ n1452 ;
  assign n1463 = n1459 & ~n1462 ;
  assign n1464 = n1463 ^ n1462 ;
  assign n1465 = ~x182 & n1458 ;
  assign n1466 = x54 & n1465 ;
  assign n1467 = n1466 ^ x180 ;
  assign n1468 = ~x180 & ~n1467 ;
  assign n1469 = ~n1464 & n1468 ;
  assign n1470 = n1469 ^ x180 ;
  assign n1471 = ~x53 & n1470 ;
  assign n1472 = x181 & ~n1471 ;
  assign n1473 = x182 & ~n487 ;
  assign n1474 = n340 & n1473 ;
  assign n1475 = n1464 & n1474 ;
  assign n1476 = n1475 ^ n1473 ;
  assign n1477 = n1476 ^ x182 ;
  assign n1478 = x183 & ~n490 ;
  assign n1479 = n341 & n1478 ;
  assign n1480 = n1462 & n1479 ;
  assign n1481 = n1480 ^ n1478 ;
  assign n1482 = n1481 ^ x183 ;
  assign n1487 = n494 & n1452 ;
  assign n1488 = n1487 ^ n493 ;
  assign n1489 = x184 & n1488 ;
  assign n1490 = n346 & n1394 ;
  assign n1491 = n323 & n1490 ;
  assign n1492 = n330 & n1491 ;
  assign n1493 = n333 & n1492 ;
  assign n1494 = ~x187 & n1493 ;
  assign n1495 = x59 & n1494 ;
  assign n1496 = x60 & n1493 ;
  assign n1497 = n514 & n1492 ;
  assign n1498 = n538 & n1491 ;
  assign n1499 = ~n731 & n1490 ;
  assign n1500 = n346 & ~n496 ;
  assign n1501 = ~n1401 & n1500 ;
  assign n1502 = n1501 ^ n496 ;
  assign n1503 = n1499 & ~n1502 ;
  assign n1504 = n1503 ^ n1502 ;
  assign n1505 = n1498 & ~n1504 ;
  assign n1506 = n1505 ^ n1504 ;
  assign n1507 = n1497 & ~n1506 ;
  assign n1508 = n1507 ^ n1506 ;
  assign n1509 = n1496 & ~n1508 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1511 = n1495 & ~n1510 ;
  assign n1512 = n1511 ^ n1510 ;
  assign n1513 = ~x186 & n1494 ;
  assign n1514 = x58 & n1513 ;
  assign n1515 = n1514 ^ x184 ;
  assign n1516 = ~x184 & ~n1515 ;
  assign n1517 = ~n1512 & n1516 ;
  assign n1518 = n1517 ^ x184 ;
  assign n1519 = ~x57 & n1518 ;
  assign n1520 = x185 & ~n1519 ;
  assign n1521 = x186 & ~n499 ;
  assign n1522 = n334 & n1521 ;
  assign n1523 = n1512 & n1522 ;
  assign n1524 = n1523 ^ n1521 ;
  assign n1525 = n1524 ^ x186 ;
  assign n1526 = x187 & ~n502 ;
  assign n1527 = n335 & n1526 ;
  assign n1528 = n1510 & n1527 ;
  assign n1529 = n1528 ^ n1526 ;
  assign n1530 = n1529 ^ x187 ;
  assign n1531 = x188 & ~n505 ;
  assign n1532 = n336 & n1531 ;
  assign n1533 = n1508 & n1532 ;
  assign n1534 = n1533 ^ n1531 ;
  assign n1535 = n1534 ^ x188 ;
  assign n1536 = n336 & ~n1506 ;
  assign n1544 = n1492 & n1536 ;
  assign n1545 = x64 & n1544 ;
  assign n1546 = n1545 ^ x64 ;
  assign n1537 = n1536 ^ n336 ;
  assign n1538 = n1537 ^ x64 ;
  assign n1547 = n1546 ^ n1538 ;
  assign n1548 = ~n505 & ~n1547 ;
  assign n1549 = ~x191 & n336 ;
  assign n1550 = n1492 & n1549 ;
  assign n1551 = x63 & n1550 ;
  assign n1552 = n1548 & n1551 ;
  assign n1553 = n1552 ^ n1548 ;
  assign n1554 = ~x190 & n1550 ;
  assign n1555 = x62 & n1554 ;
  assign n1556 = n1555 ^ x188 ;
  assign n1557 = ~x188 & ~n1556 ;
  assign n1558 = n1553 & n1557 ;
  assign n1559 = n1558 ^ x188 ;
  assign n1560 = ~x61 & n1559 ;
  assign n1561 = x189 & ~n1560 ;
  assign n1562 = x190 & ~n508 ;
  assign n1563 = n331 & n1562 ;
  assign n1564 = ~n1553 & n1563 ;
  assign n1565 = n1564 ^ n1562 ;
  assign n1566 = n1565 ^ x190 ;
  assign n1567 = x191 & ~n511 ;
  assign n1568 = n332 & n1567 ;
  assign n1569 = ~n1548 & n1568 ;
  assign n1570 = n1569 ^ n1567 ;
  assign n1571 = n1570 ^ x191 ;
  assign n1572 = x192 & ~n517 ;
  assign n1573 = n337 & n1572 ;
  assign n1574 = n1506 & n1573 ;
  assign n1575 = n1574 ^ n1572 ;
  assign n1576 = n1575 ^ x192 ;
  assign n1577 = ~x65 & x193 ;
  assign n1578 = n337 & n1491 ;
  assign n1579 = n326 & n1578 ;
  assign n1580 = x68 & n1579 ;
  assign n1581 = n535 & n1578 ;
  assign n1582 = n337 & ~n517 ;
  assign n1583 = n1504 & n1582 ;
  assign n1584 = n1583 ^ n517 ;
  assign n1585 = n1581 & ~n1584 ;
  assign n1586 = n1585 ^ n1584 ;
  assign n1587 = n1580 & ~n1586 ;
  assign n1588 = n1587 ^ n1586 ;
  assign n1589 = ~x192 & ~n1588 ;
  assign n1593 = ~x195 & n1579 ;
  assign n1594 = n1589 & n1593 ;
  assign n1597 = n521 & n1594 ;
  assign n1590 = n1589 ^ x192 ;
  assign n1598 = n1597 ^ n1590 ;
  assign n1599 = n1577 & n1598 ;
  assign n1600 = n1599 ^ x193 ;
  assign n1601 = ~x65 & ~x193 ;
  assign n1606 = x67 & n1594 ;
  assign n1607 = n1606 ^ n1590 ;
  assign n1608 = n1601 & n1607 ;
  assign n1609 = n1608 ^ x193 ;
  assign n1610 = ~x66 & n1609 ;
  assign n1611 = x194 & ~n1610 ;
  assign n1612 = x195 & ~n523 ;
  assign n1613 = n328 & n1612 ;
  assign n1614 = n1588 & n1613 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1616 = n1615 ^ x195 ;
  assign n1617 = x196 & ~n526 ;
  assign n1618 = n329 & n1617 ;
  assign n1619 = n1586 & n1618 ;
  assign n1620 = n1619 ^ n1617 ;
  assign n1621 = n1620 ^ x196 ;
  assign n1622 = ~x69 & x197 ;
  assign n1640 = ~x199 & n329 ;
  assign n1623 = n329 & ~n1584 ;
  assign n1631 = n1578 & n1623 ;
  assign n1632 = x72 & n1631 ;
  assign n1633 = n1632 ^ x72 ;
  assign n1624 = n1623 ^ n329 ;
  assign n1625 = n1624 ^ x72 ;
  assign n1634 = n1633 ^ n1625 ;
  assign n1635 = ~n526 & ~n1634 ;
  assign n1636 = ~x196 & n1635 ;
  assign n1641 = n1578 & n1636 ;
  assign n1642 = n1640 & n1641 ;
  assign n1645 = n530 & n1642 ;
  assign n1637 = n1636 ^ x196 ;
  assign n1646 = n1645 ^ n1637 ;
  assign n1647 = n1622 & n1646 ;
  assign n1648 = n1647 ^ x197 ;
  assign n1649 = ~x69 & ~x197 ;
  assign n1654 = x71 & n1642 ;
  assign n1655 = n1654 ^ n1637 ;
  assign n1656 = n1649 & n1655 ;
  assign n1657 = n1656 ^ x197 ;
  assign n1658 = ~x70 & n1657 ;
  assign n1659 = x198 & ~n1658 ;
  assign n1660 = x199 & ~n532 ;
  assign n1661 = n325 & n1660 ;
  assign n1662 = ~n1635 & n1661 ;
  assign n1663 = n1662 ^ n1660 ;
  assign n1664 = n1663 ^ x199 ;
  assign n1669 = n539 & n1584 ;
  assign n1670 = n1669 ^ n538 ;
  assign n1671 = x200 & n1670 ;
  assign n1672 = n338 & n1490 ;
  assign n1673 = ~x220 & n302 ;
  assign n1674 = n1672 & n1673 ;
  assign n1675 = n602 & n1674 ;
  assign n1676 = ~n729 & n1672 ;
  assign n1677 = n338 & ~n541 ;
  assign n1678 = n1502 & n1677 ;
  assign n1679 = n1678 ^ n541 ;
  assign n1680 = n1676 & ~n1679 ;
  assign n1681 = n1680 ^ n1679 ;
  assign n1682 = n1675 & ~n1681 ;
  assign n1683 = n1682 ^ n1681 ;
  assign n1684 = n313 & n1674 ;
  assign n1685 = ~n553 & n1684 ;
  assign n1693 = n317 & n1685 ;
  assign n1694 = x75 & n1693 ;
  assign n1695 = n1694 ^ x75 ;
  assign n1686 = n1685 ^ n1684 ;
  assign n1687 = n1686 ^ x75 ;
  assign n1696 = n1695 ^ n1687 ;
  assign n1697 = ~n1683 & ~n1696 ;
  assign n1698 = ~x200 & ~n1697 ;
  assign n1699 = ~x73 & ~n1698 ;
  assign n1700 = x74 & n317 ;
  assign n1701 = n318 & n1684 ;
  assign n1702 = n1700 & n1701 ;
  assign n1703 = n1699 & ~n1702 ;
  assign n1704 = x201 & ~n1703 ;
  assign n1705 = ~x74 & x202 ;
  assign n1706 = ~x201 & n1705 ;
  assign n1707 = ~n1699 & n1706 ;
  assign n1708 = n1707 ^ n1705 ;
  assign n1709 = n1708 ^ x202 ;
  assign n1710 = n319 & n1684 ;
  assign n1711 = n319 & n1683 ;
  assign n1712 = n567 & n1711 ;
  assign n1713 = n1712 ^ n567 ;
  assign n1714 = x203 & n1713 ;
  assign n1715 = n1710 & n1714 ;
  assign n1716 = n553 & n1715 ;
  assign n1717 = n1716 ^ n1714 ;
  assign n1718 = n1717 ^ x203 ;
  assign n1719 = ~n550 & n1710 ;
  assign n1727 = x77 & n1719 ;
  assign n1728 = n315 & n1727 ;
  assign n1729 = n1728 ^ n315 ;
  assign n1720 = n1719 ^ n1710 ;
  assign n1721 = n1720 ^ n315 ;
  assign n1730 = n1729 ^ n1721 ;
  assign n1731 = n1713 & ~n1730 ;
  assign n1732 = ~x203 & ~n1731 ;
  assign n1733 = ~x76 & ~n1732 ;
  assign n1734 = x204 & ~n1733 ;
  assign n1735 = n316 & n1710 ;
  assign n1736 = n316 & ~n544 ;
  assign n1737 = ~n1713 & n1736 ;
  assign n1738 = n1737 ^ n544 ;
  assign n1739 = x205 & ~n1738 ;
  assign n1740 = n1735 & n1739 ;
  assign n1741 = n550 & n1740 ;
  assign n1742 = n1741 ^ n1739 ;
  assign n1743 = n1742 ^ x205 ;
  assign n1744 = x80 & n1735 ;
  assign n1745 = ~n1738 & n1744 ;
  assign n1746 = n1745 ^ n1738 ;
  assign n1747 = ~x207 & n1735 ;
  assign n1748 = x79 & n1747 ;
  assign n1749 = n1748 ^ x205 ;
  assign n1750 = ~x205 & ~n1749 ;
  assign n1751 = ~n1746 & n1750 ;
  assign n1752 = n1751 ^ x205 ;
  assign n1753 = ~x78 & n1752 ;
  assign n1754 = x206 & ~n1753 ;
  assign n1755 = x207 & ~n547 ;
  assign n1756 = n314 & n1755 ;
  assign n1757 = n1746 & n1756 ;
  assign n1758 = n1757 ^ n1755 ;
  assign n1759 = n1758 ^ x207 ;
  assign n1764 = n551 & n1738 ;
  assign n1765 = n1764 ^ n550 ;
  assign n1766 = x208 & n1765 ;
  assign n1767 = ~x81 & x209 ;
  assign n1793 = ~x211 & n308 ;
  assign n1768 = n320 & n1674 ;
  assign n1775 = n305 & n1768 ;
  assign n1769 = n599 & n1768 ;
  assign n1770 = n320 & ~n569 ;
  assign n1771 = n1681 & n1770 ;
  assign n1772 = n1771 ^ n569 ;
  assign n1773 = n1769 & ~n1772 ;
  assign n1774 = n1773 ^ n1772 ;
  assign n1776 = ~n587 & n1775 ;
  assign n1784 = n308 & n1776 ;
  assign n1785 = x84 & n1784 ;
  assign n1786 = n1785 ^ x84 ;
  assign n1777 = n1776 ^ n1775 ;
  assign n1778 = n1777 ^ x84 ;
  assign n1787 = n1786 ^ n1778 ;
  assign n1788 = ~n1774 & ~n1787 ;
  assign n1789 = ~x208 & n1788 ;
  assign n1794 = n1775 & n1789 ;
  assign n1795 = n1793 & n1794 ;
  assign n1798 = n573 & n1795 ;
  assign n1790 = n1789 ^ x208 ;
  assign n1799 = n1798 ^ n1790 ;
  assign n1800 = n1767 & n1799 ;
  assign n1801 = n1800 ^ x209 ;
  assign n1802 = ~x81 & ~x209 ;
  assign n1807 = x83 & n1795 ;
  assign n1808 = n1807 ^ n1790 ;
  assign n1809 = n1802 & n1808 ;
  assign n1810 = n1809 ^ x209 ;
  assign n1811 = ~x82 & n1810 ;
  assign n1812 = x210 & ~n1811 ;
  assign n1813 = x211 & ~n575 ;
  assign n1814 = n310 & n1813 ;
  assign n1815 = ~n1788 & n1814 ;
  assign n1816 = n1815 ^ n1813 ;
  assign n1817 = n1816 ^ x211 ;
  assign n1818 = n311 & n1775 ;
  assign n1819 = n311 & ~n578 ;
  assign n1820 = n1774 & n1819 ;
  assign n1821 = n1820 ^ n578 ;
  assign n1822 = x212 & ~n1821 ;
  assign n1823 = n1818 & n1822 ;
  assign n1824 = n587 & n1823 ;
  assign n1825 = n1824 ^ n1822 ;
  assign n1826 = n1825 ^ x212 ;
  assign n1827 = ~x215 & n1818 ;
  assign n1828 = x87 & n1827 ;
  assign n1829 = x88 & n1818 ;
  assign n1830 = ~n1821 & n1829 ;
  assign n1831 = n1830 ^ n1821 ;
  assign n1832 = n1828 & ~n1831 ;
  assign n1833 = n1832 ^ n1831 ;
  assign n1834 = ~x214 & n1827 ;
  assign n1835 = x86 & n1834 ;
  assign n1836 = n1835 ^ x212 ;
  assign n1837 = ~x212 & ~n1836 ;
  assign n1838 = ~n1833 & n1837 ;
  assign n1839 = n1838 ^ x212 ;
  assign n1840 = ~x85 & n1839 ;
  assign n1841 = x213 & ~n1840 ;
  assign n1842 = x214 & ~n581 ;
  assign n1843 = n306 & n1842 ;
  assign n1844 = n1833 & n1843 ;
  assign n1845 = n1844 ^ n1842 ;
  assign n1846 = n1845 ^ x214 ;
  assign n1847 = x215 & ~n584 ;
  assign n1848 = n307 & n1847 ;
  assign n1849 = n1831 & n1848 ;
  assign n1850 = n1849 ^ n1847 ;
  assign n1851 = n1850 ^ x215 ;
  assign n1856 = n588 & n1821 ;
  assign n1857 = n1856 ^ n587 ;
  assign n1858 = x216 & n1857 ;
  assign n1859 = n312 & ~n1772 ;
  assign n1867 = n1768 & n1859 ;
  assign n1868 = x92 & n1867 ;
  assign n1869 = n1868 ^ x92 ;
  assign n1860 = n1859 ^ n312 ;
  assign n1861 = n1860 ^ x92 ;
  assign n1870 = n1869 ^ n1861 ;
  assign n1871 = ~n590 & ~n1870 ;
  assign n1872 = ~x219 & n312 ;
  assign n1873 = n1768 & n1872 ;
  assign n1874 = x91 & n1873 ;
  assign n1875 = n1871 & n1874 ;
  assign n1876 = n1875 ^ n1871 ;
  assign n1877 = ~x218 & n1873 ;
  assign n1878 = x90 & n1877 ;
  assign n1879 = n1878 ^ x216 ;
  assign n1880 = ~x216 & ~n1879 ;
  assign n1881 = n1876 & n1880 ;
  assign n1882 = n1881 ^ x216 ;
  assign n1883 = ~x89 & n1882 ;
  assign n1884 = x217 & ~n1883 ;
  assign n1885 = x218 & ~n593 ;
  assign n1886 = n303 & n1885 ;
  assign n1887 = ~n1876 & n1886 ;
  assign n1888 = n1887 ^ n1885 ;
  assign n1889 = n1888 ^ x218 ;
  assign n1890 = x219 & ~n596 ;
  assign n1891 = n304 & n1890 ;
  assign n1892 = ~n1871 & n1891 ;
  assign n1893 = n1892 ^ n1890 ;
  assign n1894 = n1893 ^ x219 ;
  assign n1895 = x220 & ~n605 ;
  assign n1896 = n321 & n1895 ;
  assign n1897 = n1681 & n1896 ;
  assign n1898 = n1897 ^ n1895 ;
  assign n1899 = n1898 ^ x220 ;
  assign n1900 = ~x93 & ~n606 ;
  assign n1901 = n322 & n1679 ;
  assign n1902 = n1900 & n1901 ;
  assign n1903 = n1902 ^ n1900 ;
  assign n1904 = n322 & n1672 ;
  assign n1905 = n298 & n613 ;
  assign n1906 = n718 & n1905 ;
  assign n1907 = n1906 ^ n718 ;
  assign n1908 = n1904 & n1907 ;
  assign n1916 = n301 & n1908 ;
  assign n1917 = x95 & n1916 ;
  assign n1918 = n1917 ^ x95 ;
  assign n1909 = n1908 ^ n1904 ;
  assign n1910 = n1909 ^ x95 ;
  assign n1919 = n1918 ^ n1910 ;
  assign n1920 = n1903 & ~n1919 ;
  assign n1921 = n720 & n1904 ;
  assign n1922 = n301 & n1921 ;
  assign n1923 = n1922 ^ x221 ;
  assign n1924 = x221 & n1923 ;
  assign n1925 = n1920 & n1924 ;
  assign n1926 = n1925 ^ x221 ;
  assign n1927 = ~x94 & x222 ;
  assign n1928 = ~x221 & n1927 ;
  assign n1929 = ~n1920 & n1928 ;
  assign n1930 = n1929 ^ n1927 ;
  assign n1931 = n1930 ^ x222 ;
  assign n1932 = n273 & n1904 ;
  assign n1933 = n273 & ~n1903 ;
  assign n1934 = n721 & ~n1933 ;
  assign n1935 = x223 & n1934 ;
  assign n1936 = n1932 & n1935 ;
  assign n1937 = ~n1907 & n1936 ;
  assign n1938 = n1937 ^ n1935 ;
  assign n1939 = n1938 ^ x223 ;
  assign n1940 = ~x96 & x224 ;
  assign n1941 = ~n718 & n1932 ;
  assign n1942 = ~x223 & n1934 ;
  assign n1943 = ~n1941 & n1942 ;
  assign n1947 = n298 & n1932 ;
  assign n1948 = n1943 & n1947 ;
  assign n1951 = n611 & n1948 ;
  assign n1944 = n1943 ^ x223 ;
  assign n1952 = n1951 ^ n1944 ;
  assign n1953 = n1940 & n1952 ;
  assign n1954 = n1953 ^ x224 ;
  assign n1955 = ~x96 & ~x224 ;
  assign n1960 = x98 & n1948 ;
  assign n1961 = n1960 ^ n1944 ;
  assign n1962 = n1955 & n1961 ;
  assign n1963 = n1962 ^ x224 ;
  assign n1964 = ~x97 & n1963 ;
  assign n1965 = x225 & ~n1964 ;
  assign n1966 = n726 & ~n1933 ;
  assign n1967 = x226 & ~n614 ;
  assign n1968 = ~n1941 & n1967 ;
  assign n1969 = n1966 & n1968 ;
  assign n1970 = n1969 ^ n1967 ;
  assign n1971 = n300 & n1932 ;
  assign n1972 = n286 & n1971 ;
  assign n1973 = n288 & n1972 ;
  assign n1974 = ~x234 & n1973 ;
  assign n1975 = n294 & n1974 ;
  assign n1976 = ~n620 & n1972 ;
  assign n1977 = ~n614 & ~n1966 ;
  assign n1978 = n715 & n1971 ;
  assign n1986 = x110 & n1978 ;
  assign n1987 = n286 & n1986 ;
  assign n1988 = n1987 ^ n286 ;
  assign n1979 = n1978 ^ n1971 ;
  assign n1980 = n1979 ^ n286 ;
  assign n1989 = n1988 ^ n1980 ;
  assign n1990 = ~n1977 & ~n1989 ;
  assign n1991 = ~n1976 & n1990 ;
  assign n1992 = x107 & n1973 ;
  assign n1993 = n1991 & n1992 ;
  assign n1994 = n1993 ^ n1991 ;
  assign n1995 = ~x226 & n1994 ;
  assign n2003 = n1974 & n1995 ;
  assign n2004 = x106 & n2003 ;
  assign n2005 = n2004 ^ x106 ;
  assign n1996 = n1995 ^ x226 ;
  assign n1997 = n1996 ^ x106 ;
  assign n2006 = n2005 ^ n1997 ;
  assign n2007 = ~x99 & n2006 ;
  assign n2008 = x227 & n2007 ;
  assign n2009 = ~n644 & n2008 ;
  assign n2010 = n1975 & n2009 ;
  assign n2011 = n2010 ^ n2008 ;
  assign n2012 = n2011 ^ x227 ;
  assign n2013 = ~x105 & ~x232 ;
  assign n2018 = n626 & n629 ;
  assign n2019 = n2018 ^ x104 ;
  assign n2020 = n2013 & n2019 ;
  assign n2021 = n2020 ^ x105 ;
  assign n2022 = n1975 & n2021 ;
  assign n2023 = n2007 & ~n2022 ;
  assign n2024 = ~x227 & ~n2023 ;
  assign n2025 = ~x100 & ~n2024 ;
  assign n2026 = n631 & n1975 ;
  assign n2027 = n292 & n2026 ;
  assign n2028 = n2027 ^ x228 ;
  assign n2029 = x228 & n2028 ;
  assign n2030 = n2025 & n2029 ;
  assign n2031 = n2030 ^ x228 ;
  assign n2032 = ~x101 & ~x228 ;
  assign n2033 = ~n2025 & n2032 ;
  assign n2034 = n2033 ^ x101 ;
  assign n2035 = ~x229 & n2034 ;
  assign n2036 = n2035 ^ n2034 ;
  assign n2037 = ~x102 & x230 ;
  assign n2038 = ~n2035 & n2037 ;
  assign n2039 = n2038 ^ x230 ;
  assign n2040 = n290 & ~n628 ;
  assign n2041 = ~n2025 & n2040 ;
  assign n2042 = n2041 ^ n628 ;
  assign n2043 = ~x231 & n2042 ;
  assign n2044 = n2043 ^ n2042 ;
  assign n2045 = ~x104 & x232 ;
  assign n2046 = ~n2043 & n2045 ;
  assign n2047 = n2046 ^ x232 ;
  assign n2048 = x233 & n644 ;
  assign n2049 = n293 & n2048 ;
  assign n2050 = ~n2007 & n2049 ;
  assign n2051 = n2050 ^ n2048 ;
  assign n2052 = n2051 ^ x233 ;
  assign n2053 = x234 & n657 ;
  assign n2054 = ~n1994 & n2053 ;
  assign n2055 = n295 & n2054 ;
  assign n2056 = n2055 ^ n2053 ;
  assign n2057 = n2056 ^ x234 ;
  assign n2058 = n296 & ~n659 ;
  assign n2059 = ~n1990 & n2058 ;
  assign n2060 = n2059 ^ n659 ;
  assign n2061 = x235 & ~n2060 ;
  assign n2062 = n1976 & n2061 ;
  assign n2063 = n296 & n2062 ;
  assign n2064 = n2063 ^ n2061 ;
  assign n2065 = n2064 ^ x235 ;
  assign n2066 = ~x108 & ~x235 ;
  assign n2067 = n2060 & n2066 ;
  assign n2068 = n2067 ^ x108 ;
  assign n2069 = x109 & n287 ;
  assign n2070 = n296 & n1972 ;
  assign n2071 = n2069 & n2070 ;
  assign n2072 = ~n2068 & ~n2071 ;
  assign n2073 = x236 & ~n2072 ;
  assign n2074 = ~x109 & x237 ;
  assign n2075 = ~x236 & n2074 ;
  assign n2076 = n2068 & n2075 ;
  assign n2077 = n2076 ^ n2074 ;
  assign n2078 = n2077 ^ x237 ;
  assign n2079 = n297 & n662 ;
  assign n2080 = ~n1990 & n2079 ;
  assign n2081 = n2080 ^ n662 ;
  assign n2082 = ~x238 & ~n2081 ;
  assign n2083 = n2082 ^ n2081 ;
  assign n2084 = ~x111 & x239 ;
  assign n2085 = ~n2082 & n2084 ;
  assign n2086 = n2085 ^ x239 ;
  assign n2087 = n285 & n297 ;
  assign n2088 = n1971 & n2087 ;
  assign n2089 = n665 ^ n297 ;
  assign n2090 = n2089 ^ n285 ;
  assign n2091 = n662 ^ n297 ;
  assign n2092 = n2091 ^ n285 ;
  assign n2093 = n1977 ^ n662 ;
  assign n2094 = n2093 ^ n665 ;
  assign n2095 = n2092 & ~n2094 ;
  assign n2096 = ~n2090 & n2095 ;
  assign n2097 = n2096 ^ n662 ;
  assign n2098 = n2097 ^ n665 ;
  assign n2099 = n285 & ~n2098 ;
  assign n2100 = ~n665 & n2099 ;
  assign n2101 = n2100 ^ n665 ;
  assign n2102 = x240 & ~n2101 ;
  assign n2103 = n2088 & n2102 ;
  assign n2104 = ~n712 & n2103 ;
  assign n2105 = n2104 ^ n2102 ;
  assign n2106 = n2105 ^ x240 ;
  assign n2107 = ~x113 & x241 ;
  assign n2108 = ~n709 & n2088 ;
  assign n2109 = ~n2101 & n2108 ;
  assign n2110 = n2109 ^ n2101 ;
  assign n2111 = n279 & n2088 ;
  assign n2112 = x117 & n2111 ;
  assign n2113 = ~n2110 & n2112 ;
  assign n2114 = n2113 ^ n2110 ;
  assign n2115 = ~x244 & n2111 ;
  assign n2116 = x116 & n2115 ;
  assign n2117 = ~n2114 & n2116 ;
  assign n2118 = n2117 ^ n2114 ;
  assign n2119 = ~x240 & ~n2118 ;
  assign n2123 = ~x243 & n2115 ;
  assign n2124 = n2119 & n2123 ;
  assign n2127 = n669 & n2124 ;
  assign n2120 = n2119 ^ x240 ;
  assign n2128 = n2127 ^ n2120 ;
  assign n2129 = n2107 & n2128 ;
  assign n2130 = n2129 ^ x241 ;
  assign n2131 = ~x113 & ~x241 ;
  assign n2136 = x115 & n2124 ;
  assign n2137 = n2136 ^ n2120 ;
  assign n2138 = n2131 & n2137 ;
  assign n2139 = n2138 ^ x241 ;
  assign n2140 = ~x114 & n2139 ;
  assign n2141 = x242 & ~n2140 ;
  assign n2142 = x243 & ~n671 ;
  assign n2143 = n281 & n2142 ;
  assign n2144 = n2118 & n2143 ;
  assign n2145 = n2144 ^ n2142 ;
  assign n2146 = n2145 ^ x243 ;
  assign n2147 = x244 & ~n674 ;
  assign n2148 = n282 & n2147 ;
  assign n2149 = n2114 & n2148 ;
  assign n2150 = n2149 ^ n2147 ;
  assign n2151 = n2150 ^ x244 ;
  assign n2152 = x245 & ~n677 ;
  assign n2153 = n283 & n2152 ;
  assign n2154 = n2110 & n2153 ;
  assign n2155 = n2154 ^ n2152 ;
  assign n2156 = n2155 ^ x245 ;
  assign n2157 = ~x245 & n283 ;
  assign n2158 = n2088 & n2157 ;
  assign n2159 = n283 ^ x245 ;
  assign n2160 = n2159 ^ x118 ;
  assign n2161 = n677 ^ n283 ;
  assign n2162 = n2161 ^ x118 ;
  assign n2163 = n2101 ^ n677 ;
  assign n2164 = n2163 ^ x245 ;
  assign n2165 = n2162 & n2164 ;
  assign n2166 = n2160 & n2165 ;
  assign n2167 = n2166 ^ n677 ;
  assign n2168 = n2167 ^ x245 ;
  assign n2169 = ~x118 & n2168 ;
  assign n2170 = ~x245 & n2169 ;
  assign n2171 = n2170 ^ x118 ;
  assign n2172 = x246 & ~n2171 ;
  assign n2173 = n2158 & n2172 ;
  assign n2174 = ~n707 & n2173 ;
  assign n2175 = n2174 ^ n2172 ;
  assign n2176 = n2175 ^ x246 ;
  assign n2177 = ~x246 & n2158 ;
  assign n2178 = ~x119 & ~x246 ;
  assign n2179 = n2171 & n2178 ;
  assign n2180 = n2179 ^ x119 ;
  assign n2181 = x247 & ~n2180 ;
  assign n2182 = n2177 & n2181 ;
  assign n2183 = ~n704 & n2182 ;
  assign n2184 = n2183 ^ n2181 ;
  assign n2185 = n2184 ^ x247 ;
  assign n2186 = n276 & n2177 ;
  assign n2187 = ~x247 & ~n2180 ;
  assign n2195 = n2177 & n2187 ;
  assign n2196 = x124 & n2195 ;
  assign n2197 = n2196 ^ x124 ;
  assign n2188 = n2187 ^ x247 ;
  assign n2189 = n2188 ^ x124 ;
  assign n2198 = n2197 ^ n2189 ;
  assign n2199 = ~x120 & n2198 ;
  assign n2200 = x248 & n2199 ;
  assign n2201 = ~n691 & n2200 ;
  assign n2202 = n2186 & n2201 ;
  assign n2203 = n2202 ^ n2200 ;
  assign n2204 = n2203 ^ x248 ;
  assign n2205 = ~x248 & n2199 ;
  assign n2213 = n2186 & n2205 ;
  assign n2214 = x123 & n2213 ;
  assign n2215 = n2214 ^ x123 ;
  assign n2206 = n2205 ^ x248 ;
  assign n2207 = n2206 ^ x123 ;
  assign n2216 = n2215 ^ n2207 ;
  assign n2217 = ~x121 & n2216 ;
  assign n2218 = n274 & n2186 ;
  assign n2219 = x122 & n2218 ;
  assign n2220 = n2219 ^ x249 ;
  assign n2221 = x249 & n2220 ;
  assign n2222 = n2217 & n2221 ;
  assign n2223 = n2222 ^ x249 ;
  assign n2224 = ~x122 & x250 ;
  assign n2225 = ~x249 & n2224 ;
  assign n2226 = ~n2217 & n2225 ;
  assign n2227 = n2226 ^ n2224 ;
  assign n2228 = n2227 ^ x250 ;
  assign n2229 = x251 & n691 ;
  assign n2230 = n275 & n2229 ;
  assign n2231 = ~n2199 & n2230 ;
  assign n2232 = n2231 ^ n2229 ;
  assign n2233 = n2232 ^ x251 ;
  assign n2234 = n347 & n737 ;
  assign n2235 = n1502 & n2234 ;
  assign n2236 = n2235 ^ n737 ;
  assign n2237 = ~x252 & ~n2236 ;
  assign n2238 = n2237 ^ n2236 ;
  assign n2239 = ~x125 & x253 ;
  assign n2240 = ~n2237 & n2239 ;
  assign n2241 = n2240 ^ x253 ;
  assign n2242 = n347 & n1399 ;
  assign n2250 = n1393 & n2242 ;
  assign n2251 = x127 & n2250 ;
  assign n2252 = n2251 ^ x127 ;
  assign n2243 = n2242 ^ n347 ;
  assign n2244 = n2243 ^ x127 ;
  assign n2253 = n2252 ^ n2244 ;
  assign n2254 = n737 & ~n2253 ;
  assign n2255 = n271 & ~n2254 ;
  assign n2256 = ~n740 & ~n2255 ;
  assign n2257 = x254 & ~n2256 ;
  assign n2262 = n747 & ~n1399 ;
  assign n2263 = n2262 ^ n746 ;
  assign n2264 = x255 & n2263 ;
  assign n2265 = n348 & n1393 ;
  assign y0 = n841 ;
  assign y1 = n853 ;
  assign y2 = n873 ;
  assign y3 = n879 ;
  assign y4 = n895 ;
  assign y5 = n901 ;
  assign y6 = ~n904 ;
  assign y7 = ~n907 ;
  assign y8 = n910 ;
  assign y9 = n915 ;
  assign y10 = n934 ;
  assign y11 = n957 ;
  assign y12 = n962 ;
  assign y13 = n971 ;
  assign y14 = n991 ;
  assign y15 = n1014 ;
  assign y16 = n1019 ;
  assign y17 = n1024 ;
  assign y18 = n1029 ;
  assign y19 = n1058 ;
  assign y20 = n1063 ;
  assign y21 = n1073 ;
  assign y22 = n1087 ;
  assign y23 = n1097 ;
  assign y24 = n1102 ;
  assign y25 = n1111 ;
  assign y26 = n1120 ;
  assign y27 = n1136 ;
  assign y28 = n1145 ;
  assign y29 = n1172 ;
  assign y30 = n1183 ;
  assign y31 = n1188 ;
  assign y32 = n1197 ;
  assign y33 = n1224 ;
  assign y34 = n1235 ;
  assign y35 = n1240 ;
  assign y36 = n1249 ;
  assign y37 = n1276 ;
  assign y38 = n1287 ;
  assign y39 = n1292 ;
  assign y40 = n1301 ;
  assign y41 = n1321 ;
  assign y42 = n1330 ;
  assign y43 = n1349 ;
  assign y44 = n1358 ;
  assign y45 = n1372 ;
  assign y46 = n1382 ;
  assign y47 = n1387 ;
  assign y48 = n1392 ;
  assign y49 = n1438 ;
  assign y50 = n1443 ;
  assign y51 = n1448 ;
  assign y52 = n1457 ;
  assign y53 = n1472 ;
  assign y54 = n1477 ;
  assign y55 = n1482 ;
  assign y56 = n1489 ;
  assign y57 = n1520 ;
  assign y58 = n1525 ;
  assign y59 = n1530 ;
  assign y60 = n1535 ;
  assign y61 = n1561 ;
  assign y62 = n1566 ;
  assign y63 = n1571 ;
  assign y64 = n1576 ;
  assign y65 = n1600 ;
  assign y66 = n1611 ;
  assign y67 = n1616 ;
  assign y68 = n1621 ;
  assign y69 = n1648 ;
  assign y70 = n1659 ;
  assign y71 = n1664 ;
  assign y72 = n1671 ;
  assign y73 = n1704 ;
  assign y74 = n1709 ;
  assign y75 = n1718 ;
  assign y76 = n1734 ;
  assign y77 = n1743 ;
  assign y78 = n1754 ;
  assign y79 = n1759 ;
  assign y80 = n1766 ;
  assign y81 = n1801 ;
  assign y82 = n1812 ;
  assign y83 = n1817 ;
  assign y84 = n1826 ;
  assign y85 = n1841 ;
  assign y86 = n1846 ;
  assign y87 = n1851 ;
  assign y88 = n1858 ;
  assign y89 = n1884 ;
  assign y90 = n1889 ;
  assign y91 = n1894 ;
  assign y92 = n1899 ;
  assign y93 = n1926 ;
  assign y94 = n1931 ;
  assign y95 = n1939 ;
  assign y96 = n1954 ;
  assign y97 = n1965 ;
  assign y98 = n1970 ;
  assign y99 = n2012 ;
  assign y100 = n2031 ;
  assign y101 = n2036 ;
  assign y102 = n2039 ;
  assign y103 = n2044 ;
  assign y104 = n2047 ;
  assign y105 = n2052 ;
  assign y106 = n2057 ;
  assign y107 = n2065 ;
  assign y108 = n2073 ;
  assign y109 = n2078 ;
  assign y110 = ~n2083 ;
  assign y111 = n2086 ;
  assign y112 = n2106 ;
  assign y113 = n2130 ;
  assign y114 = n2141 ;
  assign y115 = n2146 ;
  assign y116 = n2151 ;
  assign y117 = n2156 ;
  assign y118 = n2176 ;
  assign y119 = n2185 ;
  assign y120 = n2204 ;
  assign y121 = n2223 ;
  assign y122 = n2228 ;
  assign y123 = n2233 ;
  assign y124 = ~n2238 ;
  assign y125 = n2241 ;
  assign y126 = n2257 ;
  assign y127 = n2264 ;
  assign y128 = ~n2265 ;
endmodule
