module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n209 , n210 , n211 , n212 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 ;
  assign n65 = x21 & ~x53 ;
  assign n67 = ~x22 & x54 ;
  assign n66 = x54 ^ x22 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = ~n65 & ~n68 ;
  assign n70 = x23 & ~x55 ;
  assign n71 = n69 & n70 ;
  assign n72 = n71 ^ n69 ;
  assign n74 = x20 & ~x52 ;
  assign n73 = x52 ^ x20 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = x53 ^ x21 ;
  assign n77 = n76 ^ n65 ;
  assign n78 = ~n75 & ~n77 ;
  assign n79 = n72 & n78 ;
  assign n80 = n79 ^ n72 ;
  assign n81 = x55 ^ x23 ;
  assign n82 = n67 ^ x55 ;
  assign n83 = ~n81 & n82 ;
  assign n84 = n83 ^ x55 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = n72 & ~n74 ;
  assign n87 = x17 & ~x49 ;
  assign n89 = ~x18 & x50 ;
  assign n88 = x50 ^ x18 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = ~n87 & ~n90 ;
  assign n92 = x19 & ~x51 ;
  assign n93 = n91 & n92 ;
  assign n94 = n93 ^ n91 ;
  assign n96 = x16 & ~x48 ;
  assign n95 = x48 ^ x16 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = x49 ^ x17 ;
  assign n99 = n98 ^ n87 ;
  assign n100 = ~n97 & ~n99 ;
  assign n101 = n94 & n100 ;
  assign n102 = n101 ^ n94 ;
  assign n103 = n86 & ~n102 ;
  assign n104 = x51 ^ x19 ;
  assign n105 = n89 ^ x19 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = n106 ^ x19 ;
  assign n108 = n103 & n107 ;
  assign n109 = n108 ^ n86 ;
  assign n110 = n85 & ~n109 ;
  assign n111 = x27 & ~x59 ;
  assign n112 = x25 & x57 ;
  assign n113 = n112 ^ x25 ;
  assign n114 = ~n111 & ~n113 ;
  assign n115 = x26 & ~x58 ;
  assign n116 = n114 & n115 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = x56 & n117 ;
  assign n119 = ~x24 & n117 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = x28 & ~x60 ;
  assign n122 = ~x31 & ~n121 ;
  assign n123 = x63 & n122 ;
  assign n124 = n123 ^ x29 ;
  assign n125 = n123 ^ n121 ;
  assign n126 = ~x61 & ~n125 ;
  assign n127 = n124 & n126 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = x30 & ~x62 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = ~n120 & ~n131 ;
  assign n133 = ~n110 & n132 ;
  assign n134 = n120 ^ n118 ;
  assign n135 = n134 ^ n119 ;
  assign n136 = x59 ^ x27 ;
  assign n137 = x58 ^ x57 ;
  assign n138 = n137 ^ n111 ;
  assign n139 = n138 ^ n112 ;
  assign n142 = x59 ^ x26 ;
  assign n140 = x59 ^ x58 ;
  assign n141 = n140 ^ n111 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = ~n139 & ~n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = ~n136 & n145 ;
  assign n147 = n146 ^ x27 ;
  assign n148 = ~n131 & n147 ;
  assign n149 = n135 & n148 ;
  assign n150 = n149 ^ n131 ;
  assign n151 = ~n133 & n150 ;
  assign n152 = x63 ^ x31 ;
  assign n154 = x60 ^ x28 ;
  assign n155 = n154 ^ n121 ;
  assign n156 = n155 ^ x62 ;
  assign n153 = x62 ^ x29 ;
  assign n157 = n156 ^ n153 ;
  assign n158 = x62 ^ x61 ;
  assign n159 = n158 ^ n156 ;
  assign n160 = ~n157 & n159 ;
  assign n161 = n160 ^ n156 ;
  assign n163 = x63 ^ x30 ;
  assign n162 = x63 ^ x62 ;
  assign n164 = n163 ^ n162 ;
  assign n165 = ~n161 & ~n164 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = ~n152 & ~n166 ;
  assign n168 = n167 ^ x31 ;
  assign n169 = x45 ^ x13 ;
  assign n171 = x12 & ~x44 ;
  assign n170 = x44 ^ x12 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = n172 ^ x45 ;
  assign n174 = ~n169 & ~n173 ;
  assign n175 = n174 ^ x13 ;
  assign n176 = ~n169 & ~n171 ;
  assign n177 = x43 ^ x11 ;
  assign n179 = x42 ^ x10 ;
  assign n182 = ~x9 & x41 ;
  assign n183 = n182 ^ x43 ;
  assign n178 = x43 ^ x42 ;
  assign n184 = n183 ^ n178 ;
  assign n185 = ~n179 & n184 ;
  assign n186 = n185 ^ n178 ;
  assign n187 = ~n177 & n186 ;
  assign n188 = n187 ^ x43 ;
  assign n189 = x47 ^ x15 ;
  assign n190 = x14 & ~x46 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = ~n177 & ~n179 ;
  assign n193 = x41 ^ x9 ;
  assign n194 = n193 ^ n182 ;
  assign n197 = ~x8 & ~n194 ;
  assign n198 = n192 & n197 ;
  assign n195 = x40 & ~n194 ;
  assign n196 = n192 & n195 ;
  assign n199 = n198 ^ n196 ;
  assign n200 = x38 ^ x6 ;
  assign n201 = x7 & ~x39 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = x5 & x37 ;
  assign n204 = n203 ^ x5 ;
  assign n205 = n202 & ~n204 ;
  assign n206 = x36 ^ x4 ;
  assign n209 = x34 ^ x2 ;
  assign n211 = x34 ^ x1 ;
  assign n210 = x34 ^ x33 ;
  assign n212 = n211 ^ n210 ;
  assign n214 = x0 & ~x32 ;
  assign n215 = n214 ^ x1 ;
  assign n216 = ~n212 & n215 ;
  assign n217 = n216 ^ n211 ;
  assign n218 = ~n209 & n217 ;
  assign n207 = x35 ^ x2 ;
  assign n219 = n218 ^ n207 ;
  assign n221 = x36 ^ x3 ;
  assign n220 = x36 ^ x35 ;
  assign n222 = n221 ^ n220 ;
  assign n223 = n219 & ~n222 ;
  assign n224 = n223 ^ n221 ;
  assign n225 = ~n206 & n224 ;
  assign n226 = n225 ^ x4 ;
  assign n227 = n205 & ~n226 ;
  assign n228 = x39 ^ x7 ;
  assign n229 = n201 ^ n200 ;
  assign n232 = x39 ^ x6 ;
  assign n230 = x39 ^ x37 ;
  assign n231 = n230 ^ n203 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = ~n229 & ~n233 ;
  assign n235 = n234 ^ n232 ;
  assign n236 = ~n228 & n235 ;
  assign n237 = n236 ^ x7 ;
  assign n238 = ~n227 & n237 ;
  assign n239 = n238 ^ n196 ;
  assign n240 = n199 & n239 ;
  assign n241 = n240 ^ n198 ;
  assign n242 = n191 & ~n241 ;
  assign n243 = ~n188 & n242 ;
  assign n244 = n243 ^ n191 ;
  assign n245 = n176 & n244 ;
  assign n246 = n245 ^ n191 ;
  assign n247 = n175 & n246 ;
  assign n248 = n247 ^ n191 ;
  assign n249 = x46 ^ x14 ;
  assign n250 = n249 ^ n190 ;
  assign n251 = n250 ^ x47 ;
  assign n252 = ~n189 & ~n251 ;
  assign n253 = n252 ^ x15 ;
  assign n254 = ~n96 & n253 ;
  assign n255 = ~n248 & n254 ;
  assign n256 = n255 ^ n96 ;
  assign n257 = n94 & ~n256 ;
  assign n258 = n86 & n257 ;
  assign n259 = n132 & n258 ;
  assign n260 = ~n168 & ~n259 ;
  assign n261 = n151 & n260 ;
  assign y0 = ~n261 ;
endmodule
