module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
output y0;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, y0;
assign n_0 = x32 ^ x0;
assign n_1 = x33 ^ x1;
assign n_2 = x34 ^ x2;
assign n_3 = x35 ^ x3;
assign n_4 = x36 ^ x4;
assign n_5 = x37 ^ x5;
assign n_6 = x38 ^ x6;
assign n_7 = ~x6 & x38;
assign n_8 = x39 ^ x7;
assign n_9 = ~x7 ^ x39;
assign n_10 = x41 ^ x9;
assign n_11 = x9 & ~x41;
assign n_12 = ~x10 & x42;
assign n_13 = x42 ^ x10;
assign n_14 = ~x11 & x43;
assign n_15 = x43 ^ x11;
assign n_16 = ~x12 ^ x44;
assign n_17 = x45 ^ x13;
assign n_18 = ~x14 & x46;
assign n_19 = x46 ^ x14;
assign n_20 = ~x15 & x47;
assign n_21 = x47 ^ x15;
assign n_22 = x48 ^ x16;
assign n_23 = ~x16 & x48;
assign n_24 = x49 ^ x17;
assign n_25 = ~x17 ^ x49;
assign n_26 = ~x18 & x50;
assign n_27 = x51 ^ x19;
assign n_28 = ~x19 ^ x51;
assign n_29 = x52 ^ x20;
assign n_30 = ~x20 & x52;
assign n_31 = x53 ^ x21;
assign n_32 = ~x21 & x53;
assign n_33 = x54 ^ x22;
assign n_34 = ~x22 & x54;
assign n_35 = x55 ^ x23;
assign n_36 = ~x23 & x55;
assign n_37 = x57 ^ x25;
assign n_38 = x58 ^ x26;
assign n_39 = ~x26 & x58;
assign n_40 = x59 ^ x27;
assign n_41 = ~x27 & x59;
assign n_42 = ~x28 & x60;
assign n_43 = x60 ^ x28;
assign n_44 = ~x29 & x61;
assign n_45 = x61 ^ x29;
assign n_46 = ~x30 & x62;
assign n_47 = x31 & ~x63;
assign n_48 = x63 ^ x31;
assign n_49 = x32 & ~n_0;
assign n_50 = n_6 ^ n_7;
assign n_51 = ~n_7 & n_9;
assign n_52 = n_10 ^ n_11;
assign n_53 = n_11 ^ x42;
assign n_54 = ~n_12 & ~n_14;
assign n_55 = ~x45 & ~n_17;
assign n_56 = ~n_18 & ~n_20;
assign n_57 = n_19 ^ n_20;
assign n_58 = n_22 ^ n_23;
assign n_59 = n_26 ^ x18;
assign n_60 = ~n_26 & n_28;
assign n_61 = n_29 ^ n_30;
assign n_62 = ~n_30 & ~n_32;
assign n_63 = n_33 ^ n_34;
assign n_64 = ~n_34 & ~n_36;
assign n_65 = ~x57 & ~n_37;
assign n_66 = n_38 ^ n_41;
assign n_67 = ~n_41 & ~n_39;
assign n_68 = n_43 ^ n_42;
assign n_69 = ~n_42 & ~n_44;
assign n_70 = n_46 ^ x30;
assign n_71 = ~n_46 & ~n_47;
assign n_72 = n_49 ^ x1;
assign n_73 = n_50 ^ x39;
assign n_74 = ~x40 & ~n_52;
assign n_75 = x8 & ~n_52;
assign n_76 = ~n_13 & ~n_53;
assign n_77 = n_55 ^ x13;
assign n_78 = n_55 ^ x14;
assign n_79 = n_58 ^ x49;
assign n_80 = n_59 ^ x50;
assign n_81 = n_61 ^ x53;
assign n_82 = n_63 ^ x55;
assign n_83 = n_64 & n_62;
assign n_84 = n_65 ^ x26;
assign n_85 = n_65 ^ x25;
assign n_86 = n_68 ^ x61;
assign n_87 = n_70 ^ x62;
assign n_88 = n_69 & n_71;
assign n_89 = n_72 ^ x32;
assign n_90 = ~n_8 & n_73;
assign n_91 = n_74 & n_54;
assign n_92 = n_54 & n_75;
assign n_93 = n_76 ^ x42;
assign n_94 = n_56 & n_77;
assign n_95 = n_78 ^ x45;
assign n_96 = ~n_24 & n_79;
assign n_97 = ~n_31 & n_81;
assign n_98 = ~n_35 & n_82;
assign n_99 = n_84 ^ x57;
assign n_100 = n_67 & n_85;
assign n_101 = ~n_45 & n_86;
assign n_102 = n_1 & ~n_89;
assign n_103 = n_90 ^ x7;
assign n_104 = x8 & n_91;
assign n_105 = n_92 ^ n_91;
assign n_106 = n_93 ^ x43;
assign n_107 = x12 & n_94;
assign n_108 = n_57 & ~n_95;
assign n_109 = n_96 ^ x17;
assign n_110 = n_97 ^ x21;
assign n_111 = n_98 ^ x23;
assign n_112 = n_66 & ~n_99;
assign n_113 = ~x56 & n_100;
assign n_114 = x24 & n_100;
assign n_115 = n_101 ^ x29;
assign n_116 = n_102 ^ n_49;
assign n_117 = ~n_15 & n_106;
assign n_118 = ~x44 & n_107;
assign n_119 = n_108 ^ n_55;
assign n_120 = n_109 ^ x51;
assign n_121 = n_64 & n_110;
assign n_122 = n_112 ^ n_65;
assign n_123 = ~n_113 & ~n_114;
assign n_124 = n_115 ^ x63;
assign n_125 = n_116 ^ x32;
assign n_126 = n_117 ^ x43;
assign n_127 = n_119 ^ x45;
assign n_128 = n_120 ^ x51;
assign n_129 = n_122 ^ x57;
assign n_130 = n_123 ^ n_113;
assign n_131 = n_88 & ~n_123;
assign n_132 = n_124 ^ x63;
assign n_133 = n_125 ^ x34;
assign n_134 = ~n_104 & n_126;
assign n_135 = n_127 ^ x47;
assign n_136 = ~n_26 & n_128;
assign n_137 = n_129 ^ x59;
assign n_138 = n_130 ^ n_114;
assign n_139 = ~n_46 & n_132;
assign n_140 = ~n_2 & n_133;
assign n_141 = ~n_21 & n_135;
assign n_142 = n_136 ^ x50;
assign n_143 = n_136 ^ x51;
assign n_144 = ~n_40 & n_137;
assign n_145 = n_139 ^ x62;
assign n_146 = n_139 ^ x63;
assign n_147 = n_140 ^ x34;
assign n_148 = n_141 ^ x47;
assign n_149 = n_142 & n_80;
assign n_150 = n_144 ^ x59;
assign n_151 = n_145 & n_87;
assign n_152 = n_147 ^ x35;
assign n_153 = ~n_118 & n_148;
assign n_154 = n_149 ^ n_59;
assign n_155 = n_150 & n_138;
assign n_156 = n_151 ^ n_70;
assign n_157 = ~n_3 & n_152;
assign n_158 = n_154 ^ n_143;
assign n_159 = n_88 & ~n_155;
assign n_160 = n_156 ^ n_146;
assign n_161 = n_157 ^ x35;
assign n_162 = n_158 ^ x50;
assign n_163 = n_160 ^ x62;
assign n_164 = n_161 ^ x36;
assign n_165 = ~n_27 & n_162;
assign n_166 = ~n_48 & ~n_163;
assign n_167 = ~n_4 & n_164;
assign n_168 = n_165 ^ x19;
assign n_169 = n_166 ^ x31;
assign n_170 = n_167 ^ x36;
assign n_171 = n_83 & n_168;
assign n_172 = n_170 ^ x37;
assign n_173 = ~n_121 & ~n_171;
assign n_174 = ~n_5 & n_172;
assign n_175 = ~n_111 & n_173;
assign n_176 = n_174 ^ x37;
assign n_177 = n_131 & ~n_175;
assign n_178 = n_51 & ~n_176;
assign n_179 = ~n_159 & ~n_177;
assign n_180 = ~n_103 & ~n_178;
assign n_181 = n_105 & ~n_180;
assign n_182 = n_134 & ~n_181;
assign n_183 = n_16 & ~n_182;
assign n_184 = n_94 & n_183;
assign n_185 = n_153 & ~n_184;
assign n_186 = ~n_23 & ~n_185;
assign n_187 = n_60 & n_186;
assign n_188 = n_25 & n_187;
assign n_189 = n_83 & n_188;
assign n_190 = n_131 & n_189;
assign n_191 = n_169 & ~n_190;
assign n_192 = n_179 & n_191;
assign y0 = n_192;
endmodule